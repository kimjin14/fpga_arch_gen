//testbench for fpga_top.v
`timescale 1 ns / 1 ps

module fpga_top_tb ();

localparam N_INPUTS = 1000;
localparam SEED = 32'hBAADF00D;

	reg [7777:0]bitstream =
		7778'b10010000000010000101101001111000000000010101000001011011010001000100010000000000000000000000000000000000000000000000000010000000000000000010110110100100110011001000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101000101100110111011101100010001000100000001000000010001000100010001000000010001000100000001101110010101010101011000000000000000000000000000000010000000000000001000000000000000001010110011001100110011010000000000000000000000000000000000000000000000000000000000000000000101010101010101010101100000000000000000000000000000000000000000000000000000000000000000101011010101010101010101000000010000000100000001000000010000000000000001000000010000000000010101100110011001100110000000100000001000000000000000000000000000000000000000000000000000000000010000101010110101011011101110100000000100010001000100010001000000000000000100000000000000010000000110001000100010001000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011011101110111011101110000000000000001000000000000000000000000000000010000000000000000010101101010001000100010100010001000100010001000000010001000100000001000100010000000100000001010110010110011001101000100000000000100000000000000000000000000000000000000000000000000001010001011001100110010001000100010001000100010001000000000001000000000000000000000000000110111001010101010101100010001000100010001000100010001000000000000000100000001000000000101011010101010101010100000000000000000000000000000000000000000000000000000000010000000001011011010000100010001010001000100010001000100010001000100010001000000010000000100000000000000000010010101101010001000100010001000000000100000000000000010000000000000001000000010000000100000000000110111001100110011001100000000000000010000000000000001000000010000000100000000000000000000101010101010101010100000000000000000100000000000000010000000000000001000000000000000000011011100101010101010110000000100000001000000010000000100010001000100010001000000000000010101101001001000100010000010001000100000001000100010000000000010001000000000000000000000001100010101010101010100000000010000000100000001000000000000000100000000000000010000000001011011010010101010101010001000100000001000100010001000100000001000000010001000100010000010110110100100110011001100010001000100010001000100010000000000000000000100010001000000000101011001100110011001100000000000000000000000000000000000000000000000001000000000000000000011000101010011001100100000000000000000000000000000000000000000000100000001000000010000110000111010100001101010001000100010001010000000000000001000000000000000100000000000000000000000000000000000110111001100110011001100000000000000010000000100000001000000010000000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101101001001000100010100010001000100010001000100010001000000010000000100000000000000001000000110101010101010101000000010000000100000000000000010000000100000000000000000000000000001010001000100010001000000000000000000000000010000000000000000000000010000000100000000000110111001010101010101000010001000100000001000000010000000100000001000000010000000100000101011010101001100110011000100010001000100010001000100010001000100010001000100010000000000010101011001100110011000000000000000000000000000000000000000000000000000000000100000000010000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111001010101010101000000000000000000000000000000000000000000000000000000000000100000101011010100010001000100000000000000000000000000000000000000000000000000000000000001000000010101100110011001100100000000000000000000000000000000000000000000000000000000100000000010101100110011001100110000000000000000000000000000000000000000000000000100000000000000000001010101100110011001100000000000000000000000000000000010000000100000001000000000000000001101010100100100010001000000000000000000000100010001000000000000000000000001000000010000000110111000100010001000100000001000000010000000000000001000000010000000000000000000000000101011010101010101010101000000010000000100000000000000010000000100000001000000010000000001011011011010101010101010001000100000001000100010001000100010001000100010001000100010000000000000001010001000100100001000000111010001110000010101010101010101010101010101111111111101010101010101010111111111111111111111111111111111111111111000101010101010111111111111111111111111111000010010001010110100000000000000001010000000000000000110101010110101010101010101010101010101010101010101010000000010110000000000000000000000000000000000000001011000010001010101111111001111111110000001010100101010100011010111100000000000101011010101010010101010101111010111101010111111101011111111111111111111110101111101011111101010101000000000000000000000010000101110000000000000000000101010110101010101010010101010000001100010101010101010101010101010101010101010100001000010101000000001110101001000000000000001010100000000000000000001010101010101010101010101111111110101010101010101010100111010100110101010101011111000010101010100101010111010101011111111111110101010111000000000000000000000000000000000000000010101010101010101010000000000011110000000000001010101010101010101010101010000000000000010011011101011111110101010101011010000000000001010101011110111111111111000010010101010101010100010101011111111101010000000000010000101001010111010101010110100100100100110101000111011010101000100011010101110101000010101010100101010101000000001100101010101010101010010110100000010001000001010110010001011010100101001010101010101101010001101101101010010011101010100100000000010011101101100111100110010000000010101001000000000010101000010101010101010101010101010110100001101111010101011010100101011001010110100001111000000101001001110100001110000111110010110100100001001010101011000001101000100110010101000000101010101111010110100101010100001001101010100010101100010000101010000001101001011000001011000000000000010111011001011000100100010100100000000011000000111000000101010101000101011000001001101100101010101001010101101010011010011001101011000000100000000000101010101000100100011111101101010011000010101100001100000101011101010101010101011101100001111111010111110111010111111101010101010011111100111111111000001010100110100100010111111111111111000000000000010101010100000101011101010101010101010101001000000101010101010101010111000111011011111101010101011111111101010101010101000011111100011011111101011010100000000001010101010101000100111111100010001001100011111111010101011101111001101001110100110101010110000110000001010100001110101010101010101010011001011010000000001001100101100110100000000110101001010011011111010110011000010101000010101000010010100010000100111000000101011000010100111011011011000101011000101010000000001000001010101001000001100110001100010010010010000000000100000101010101000001001000000000101001010010010101001010100000001101001001101100011101000101100000000001011001011010010010010001010101101010100001010001010010110110100110101001100000101010101011110100000000101010000100000010101000101001100010000000000000010001001001010000001001001001010000110110100110100010100000001010001010101010101010001010101000010101010101000010100000001000000000000110100001100000101010101001011010000101011011011011001010010001010101101010010101010111111110100000010100000101101101000000110101100101010011010110000000000000000011111110101010101000000101101111011010010101010101010101000110101010001010111111111101011101;

	reg 	clk;
	reg 	reset;
	reg 	config_clk;
	reg 	config_in;
	reg 	config_en;
	wire 	config_out;
	reg 	[7:0]io_0_1_wire_reg;
	wire 	[7:0]io_0_1_wire;
	reg 	[7:0]io_0_2_wire_reg;
	wire 	[7:0]io_0_2_wire;
	reg 	[7:0]io_0_3_wire_reg;
	wire 	[7:0]io_0_3_wire;
	reg 	[7:0]io_0_4_wire_reg;
	wire 	[7:0]io_0_4_wire;
	reg 	[7:0]io_0_5_wire_reg;
	wire 	[7:0]io_0_5_wire;
	reg 	[7:0]io_1_0_wire_reg;
	wire 	[7:0]io_1_0_wire;
	reg 	[7:0]io_1_6_wire_reg;
	wire 	[7:0]io_1_6_wire;
	reg 	[7:0]io_2_0_wire_reg;
	wire 	[7:0]io_2_0_wire;
	reg 	[7:0]io_2_6_wire_reg;
	wire 	[7:0]io_2_6_wire;
	reg 	[7:0]io_3_0_wire_reg;
	wire 	[7:0]io_3_0_wire;
	reg 	[7:0]io_3_6_wire_reg;
	wire 	[7:0]io_3_6_wire;
	reg 	[7:0]io_4_0_wire_reg;
	wire 	[7:0]io_4_0_wire;
	reg 	[7:0]io_4_6_wire_reg;
	wire 	[7:0]io_4_6_wire;
	reg 	[7:0]io_5_0_wire_reg;
	wire 	[7:0]io_5_0_wire;
	reg 	[7:0]io_5_6_wire_reg;
	wire 	[7:0]io_5_6_wire;
	reg 	[7:0]io_6_1_wire_reg;
	wire 	[7:0]io_6_1_wire;
	reg 	[7:0]io_6_2_wire_reg;
	wire 	[7:0]io_6_2_wire;
	reg 	[7:0]io_6_3_wire_reg;
	wire 	[7:0]io_6_3_wire;
	reg 	[7:0]io_6_4_wire_reg;
	wire 	[7:0]io_6_4_wire;
	reg 	[7:0]io_6_5_wire_reg;
	wire 	[7:0]io_6_5_wire;

	assign io_0_1_wire = io_0_1_wire_reg;
	assign io_0_2_wire = io_0_2_wire_reg;
	assign io_0_3_wire = io_0_3_wire_reg;
	assign io_0_4_wire = io_0_4_wire_reg;
	assign io_0_5_wire = io_0_5_wire_reg;
	assign io_1_0_wire = io_1_0_wire_reg;
	assign io_1_6_wire = io_1_6_wire_reg;
	assign io_2_0_wire = io_2_0_wire_reg;
	assign io_2_6_wire = io_2_6_wire_reg;
	assign io_3_0_wire = io_3_0_wire_reg;
	assign io_3_6_wire = io_3_6_wire_reg;
	assign io_4_0_wire = io_4_0_wire_reg;
	assign io_4_6_wire = io_4_6_wire_reg;
	assign io_5_0_wire = io_5_0_wire_reg;
	assign io_5_6_wire = io_5_6_wire_reg;
	assign io_6_1_wire = io_6_1_wire_reg;
	assign io_6_2_wire = io_6_2_wire_reg;
	assign io_6_3_wire = io_6_3_wire_reg;
	assign io_6_4_wire = io_6_4_wire_reg;
	assign io_6_5_wire = io_6_5_wire_reg;

	fpga_top dut (
		.clk(clk),
		.reset(reset),
		.config_clk(config_clk),
		.config_in(config_in),
		.config_en(config_en),
		.config_out(config_out),
		.io_0_1_wire(io_0_1_wire),
		.io_0_2_wire(io_0_2_wire),
		.io_0_3_wire(io_0_3_wire),
		.io_0_4_wire(io_0_4_wire),
		.io_0_5_wire(io_0_5_wire),
		.io_1_0_wire(io_1_0_wire),
		.io_1_6_wire(io_1_6_wire),
		.io_2_0_wire(io_2_0_wire),
		.io_2_6_wire(io_2_6_wire),
		.io_3_0_wire(io_3_0_wire),
		.io_3_6_wire(io_3_6_wire),
		.io_4_0_wire(io_4_0_wire),
		.io_4_6_wire(io_4_6_wire),
		.io_5_0_wire(io_5_0_wire),
		.io_5_6_wire(io_5_6_wire),
		.io_6_1_wire(io_6_1_wire),
		.io_6_2_wire(io_6_2_wire),
		.io_6_3_wire(io_6_3_wire),
		.io_6_4_wire(io_6_4_wire),
		.io_6_5_wire(io_6_5_wire)
	);

	always begin
		#0.5
		clk = ~clk;
		config_clk = ~config_clk;
	end

	reg [31:0] prod_rand = SEED;
	integer prod_n;

	initial begin
		reset = 0;
		config_en = 0;
		clk = 0;
		config_clk = 0;
		#10;

		reset = 1;
		config_en = 1;
		for (prod_n = 0; prod_n < 7779; prod_n = prod_n + 1) begin
			@(negedge config_clk);
			config_in = bitstream[prod_n];
		end

		config_en = 0;
		for (prod_n = 0; prod_n < N_INPUTS; prod_n = prod_n + 1) begin
			@(negedge clk);
			prod_rand = $random(prod_rand);
			io_0_1_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_0_2_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_0_3_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_0_4_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_0_5_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_1_0_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_1_6_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_2_0_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_2_6_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_3_0_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_3_6_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_4_0_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_4_6_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_5_0_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_5_6_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_6_1_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_6_2_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_6_3_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_6_4_wire_reg = prod_rand;
			prod_rand = $random(prod_rand);
			io_6_5_wire_reg = prod_rand;
		end

		$finish(0);
	end

endmodule

