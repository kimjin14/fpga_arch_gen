module fpga_top (
	input clk,
	input reset,
	inout [7:0]io_0_1_wire,
	inout [7:0]io_0_2_wire,
	inout [7:0]io_0_3_wire,
	inout [7:0]io_0_4_wire,
	inout [7:0]io_0_5_wire,
	inout [7:0]io_1_0_wire,
	inout [7:0]io_1_6_wire,
	inout [7:0]io_2_0_wire,
	inout [7:0]io_2_6_wire,
	inout [7:0]io_3_0_wire,
	inout [7:0]io_3_6_wire,
	inout [7:0]io_4_0_wire,
	inout [7:0]io_4_6_wire,
	inout [7:0]io_5_0_wire,
	inout [7:0]io_5_6_wire,
	inout [7:0]io_6_1_wire,
	inout [7:0]io_6_2_wire,
	inout [7:0]io_6_3_wire,
	inout [7:0]io_6_4_wire,
	inout [7:0]io_6_5_wire,
	input config_clk,
	input config_in,
	input config_en,
	output config_out
);

wire n24; //IPIN (0,1) #0 0
wire n25; //OPIN (0,1) #1 2313 2312 2311 2310
wire n26; //IPIN (0,1) #2 2
wire n27; //IPIN (0,1) #3 3
wire n28; //OPIN (0,1) #4 2317 2316 2315 2314
wire n29; //IPIN (0,1) #5 5
wire n30; //IPIN (0,1) #6 6
wire n31; //OPIN (0,1) #7 2321 2320 2319 2318
wire n32; //IPIN (0,1) #8 8
wire n33; //IPIN (0,1) #9 9
wire n34; //OPIN (0,1) #10 2325 2324 2323 2322
wire n35; //IPIN (0,1) #11 11
wire n36; //IPIN (0,1) #12 12
wire n37; //OPIN (0,1) #13 2329 2328 2327 2326
wire n38; //IPIN (0,1) #14 14
wire n39; //IPIN (0,1) #15 15
wire n40; //OPIN (0,1) #16 2313 2312 2311 2310
wire n41; //IPIN (0,1) #17 17
wire n42; //IPIN (0,1) #18 18
wire n43; //OPIN (0,1) #19 2317 2316 2315 2314
wire n44; //IPIN (0,1) #20 20
wire n45; //IPIN (0,1) #21 21
wire n46; //OPIN (0,1) #22 2321 2320 2319 2318
wire n47; //IPIN (0,1) #23 23
wire n72; //IPIN (0,2) #0 48
wire n73; //OPIN (0,2) #1 2333 2332 2331 2330
wire n74; //IPIN (0,2) #2 50
wire n75; //IPIN (0,2) #3 51
wire n76; //OPIN (0,2) #4 2337 2336 2335 2334
wire n77; //IPIN (0,2) #5 53
wire n78; //IPIN (0,2) #6 54
wire n79; //OPIN (0,2) #7 2341 2340 2339 2338
wire n80; //IPIN (0,2) #8 56
wire n81; //IPIN (0,2) #9 57
wire n82; //OPIN (0,2) #10 2345 2344 2343 2342
wire n83; //IPIN (0,2) #11 59
wire n84; //IPIN (0,2) #12 60
wire n85; //OPIN (0,2) #13 2349 2348 2347 2346
wire n86; //IPIN (0,2) #14 62
wire n87; //IPIN (0,2) #15 63
wire n88; //OPIN (0,2) #16 2333 2332 2331 2330
wire n89; //IPIN (0,2) #17 65
wire n90; //IPIN (0,2) #18 66
wire n91; //OPIN (0,2) #19 2337 2336 2335 2334
wire n92; //IPIN (0,2) #20 68
wire n93; //IPIN (0,2) #21 69
wire n94; //OPIN (0,2) #22 2341 2340 2339 2338
wire n95; //IPIN (0,2) #23 71
wire n120; //IPIN (0,3) #0 96
wire n121; //OPIN (0,3) #1 2353 2352 2351 2350
wire n122; //IPIN (0,3) #2 98
wire n123; //IPIN (0,3) #3 99
wire n124; //OPIN (0,3) #4 2357 2356 2355 2354
wire n125; //IPIN (0,3) #5 101
wire n126; //IPIN (0,3) #6 102
wire n127; //OPIN (0,3) #7 2361 2360 2359 2358
wire n128; //IPIN (0,3) #8 104
wire n129; //IPIN (0,3) #9 105
wire n130; //OPIN (0,3) #10 2365 2364 2363 2362
wire n131; //IPIN (0,3) #11 107
wire n132; //IPIN (0,3) #12 108
wire n133; //OPIN (0,3) #13 2369 2368 2367 2366
wire n134; //IPIN (0,3) #14 110
wire n135; //IPIN (0,3) #15 111
wire n136; //OPIN (0,3) #16 2353 2352 2351 2350
wire n137; //IPIN (0,3) #17 113
wire n138; //IPIN (0,3) #18 114
wire n139; //OPIN (0,3) #19 2357 2356 2355 2354
wire n140; //IPIN (0,3) #20 116
wire n141; //IPIN (0,3) #21 117
wire n142; //OPIN (0,3) #22 2361 2360 2359 2358
wire n143; //IPIN (0,3) #23 119
wire n168; //IPIN (0,4) #0 144
wire n169; //OPIN (0,4) #1 2373 2372 2371 2370
wire n170; //IPIN (0,4) #2 146
wire n171; //IPIN (0,4) #3 147
wire n172; //OPIN (0,4) #4 2377 2376 2375 2374
wire n173; //IPIN (0,4) #5 149
wire n174; //IPIN (0,4) #6 150
wire n175; //OPIN (0,4) #7 2381 2380 2379 2378
wire n176; //IPIN (0,4) #8 152
wire n177; //IPIN (0,4) #9 153
wire n178; //OPIN (0,4) #10 2385 2384 2383 2382
wire n179; //IPIN (0,4) #11 155
wire n180; //IPIN (0,4) #12 156
wire n181; //OPIN (0,4) #13 2389 2388 2387 2386
wire n182; //IPIN (0,4) #14 158
wire n183; //IPIN (0,4) #15 159
wire n184; //OPIN (0,4) #16 2373 2372 2371 2370
wire n185; //IPIN (0,4) #17 161
wire n186; //IPIN (0,4) #18 162
wire n187; //OPIN (0,4) #19 2377 2376 2375 2374
wire n188; //IPIN (0,4) #20 164
wire n189; //IPIN (0,4) #21 165
wire n190; //OPIN (0,4) #22 2381 2380 2379 2378
wire n191; //IPIN (0,4) #23 167
wire n216; //IPIN (0,5) #0 192
wire n217; //OPIN (0,5) #1 2393 2392 2391 2390
wire n218; //IPIN (0,5) #2 194
wire n219; //IPIN (0,5) #3 195
wire n220; //OPIN (0,5) #4 2397 2396 2395 2394
wire n221; //IPIN (0,5) #5 197
wire n222; //IPIN (0,5) #6 198
wire n223; //OPIN (0,5) #7 2401 2400 2399 2398
wire n224; //IPIN (0,5) #8 200
wire n225; //IPIN (0,5) #9 201
wire n226; //OPIN (0,5) #10 2405 2404 2403 2402
wire n227; //IPIN (0,5) #11 203
wire n228; //IPIN (0,5) #12 204
wire n229; //OPIN (0,5) #13 2409 2408 2407 2406
wire n230; //IPIN (0,5) #14 206
wire n231; //IPIN (0,5) #15 207
wire n232; //OPIN (0,5) #16 2393 2392 2391 2390
wire n233; //IPIN (0,5) #17 209
wire n234; //IPIN (0,5) #18 210
wire n235; //OPIN (0,5) #19 2397 2396 2395 2394
wire n236; //IPIN (0,5) #20 212
wire n237; //IPIN (0,5) #21 213
wire n238; //OPIN (0,5) #22 2401 2400 2399 2398
wire n239; //IPIN (0,5) #23 215
wire n264; //IPIN (1,0) #0 240
wire n265; //OPIN (1,0) #1 1713 1712 1711 1710
wire n266; //IPIN (1,0) #2 242
wire n267; //IPIN (1,0) #3 243
wire n268; //OPIN (1,0) #4 1717 1716 1715 1714
wire n269; //IPIN (1,0) #5 245
wire n270; //IPIN (1,0) #6 246
wire n271; //OPIN (1,0) #7 1721 1720 1719 1718
wire n272; //IPIN (1,0) #8 248
wire n273; //IPIN (1,0) #9 249
wire n274; //OPIN (1,0) #10 1725 1724 1723 1722
wire n275; //IPIN (1,0) #11 251
wire n276; //IPIN (1,0) #12 252
wire n277; //OPIN (1,0) #13 1729 1728 1727 1726
wire n278; //IPIN (1,0) #14 254
wire n279; //IPIN (1,0) #15 255
wire n280; //OPIN (1,0) #16 1713 1712 1711 1710
wire n281; //IPIN (1,0) #17 257
wire n282; //IPIN (1,0) #18 258
wire n283; //OPIN (1,0) #19 1717 1716 1715 1714
wire n284; //IPIN (1,0) #20 260
wire n285; //IPIN (1,0) #21 261
wire n286; //OPIN (1,0) #22 1721 1720 1719 1718
wire n287; //IPIN (1,0) #23 263
wire n303; //IPIN (1,1) #0 288
wire n304; //IPIN (1,1) #1 289
wire n305; //IPIN (1,1) #2 290
wire n306; //IPIN (1,1) #3 291
wire n307; //IPIN (1,1) #4 292
wire n308; //IPIN (1,1) #5 293
wire n309; //IPIN (1,1) #6 294
wire n310; //IPIN (1,1) #7 295
wire n311; //IPIN (1,1) #8 296
wire n312; //IPIN (1,1) #9 297
wire n313; //IPIN (1,1) #10 298
wire n314; //IPIN (1,1) #11 299
wire n315; //OPIN (1,1) #12 1813 1812 1811 1810
wire n316; //OPIN (1,1) #13 2413 2412 2411 2410
wire n317; //IPIN (1,1) #14 302
wire n333; //IPIN (1,2) #0 318
wire n334; //IPIN (1,2) #1 319
wire n335; //IPIN (1,2) #2 320
wire n336; //IPIN (1,2) #3 321
wire n337; //IPIN (1,2) #4 322
wire n338; //IPIN (1,2) #5 323
wire n339; //IPIN (1,2) #6 324
wire n340; //IPIN (1,2) #7 325
wire n341; //IPIN (1,2) #8 326
wire n342; //IPIN (1,2) #9 327
wire n343; //IPIN (1,2) #10 328
wire n344; //IPIN (1,2) #11 329
wire n345; //OPIN (1,2) #12 1913 1912 1911 1910
wire n346; //OPIN (1,2) #13 2433 2432 2431 2430
wire n347; //IPIN (1,2) #14 332
wire n363; //IPIN (1,3) #0 348
wire n364; //IPIN (1,3) #1 349
wire n365; //IPIN (1,3) #2 350
wire n366; //IPIN (1,3) #3 351
wire n367; //IPIN (1,3) #4 352
wire n368; //IPIN (1,3) #5 353
wire n369; //IPIN (1,3) #6 354
wire n370; //IPIN (1,3) #7 355
wire n371; //IPIN (1,3) #8 356
wire n372; //IPIN (1,3) #9 357
wire n373; //IPIN (1,3) #10 358
wire n374; //IPIN (1,3) #11 359
wire n375; //OPIN (1,3) #12 2013 2012 2011 2010
wire n376; //OPIN (1,3) #13 2453 2452 2451 2450
wire n377; //IPIN (1,3) #14 362
wire n393; //IPIN (1,4) #0 378
wire n394; //IPIN (1,4) #1 379
wire n395; //IPIN (1,4) #2 380
wire n396; //IPIN (1,4) #3 381
wire n397; //IPIN (1,4) #4 382
wire n398; //IPIN (1,4) #5 383
wire n399; //IPIN (1,4) #6 384
wire n400; //IPIN (1,4) #7 385
wire n401; //IPIN (1,4) #8 386
wire n402; //IPIN (1,4) #9 387
wire n403; //IPIN (1,4) #10 388
wire n404; //IPIN (1,4) #11 389
wire n405; //OPIN (1,4) #12 2113 2112 2111 2110
wire n406; //OPIN (1,4) #13 2473 2472 2471 2470
wire n407; //IPIN (1,4) #14 392
wire n423; //IPIN (1,5) #0 408
wire n424; //IPIN (1,5) #1 409
wire n425; //IPIN (1,5) #2 410
wire n426; //IPIN (1,5) #3 411
wire n427; //IPIN (1,5) #4 412
wire n428; //IPIN (1,5) #5 413
wire n429; //IPIN (1,5) #6 414
wire n430; //IPIN (1,5) #7 415
wire n431; //IPIN (1,5) #8 416
wire n432; //IPIN (1,5) #9 417
wire n433; //IPIN (1,5) #10 418
wire n434; //IPIN (1,5) #11 419
wire n435; //OPIN (1,5) #12 2213 2212 2211 2210
wire n436; //OPIN (1,5) #13 2493 2492 2491 2490
wire n437; //IPIN (1,5) #14 422
wire n462; //IPIN (1,6) #0 438
wire n463; //OPIN (1,6) #1 2217 2216 2215 2214
wire n464; //IPIN (1,6) #2 440
wire n465; //IPIN (1,6) #3 441
wire n466; //OPIN (1,6) #4 2221 2220 2219 2218
wire n467; //IPIN (1,6) #5 443
wire n468; //IPIN (1,6) #6 444
wire n469; //OPIN (1,6) #7 2225 2224 2223 2222
wire n470; //IPIN (1,6) #8 446
wire n471; //IPIN (1,6) #9 447
wire n472; //OPIN (1,6) #10 2229 2228 2227 2226
wire n473; //IPIN (1,6) #11 449
wire n474; //IPIN (1,6) #12 450
wire n475; //OPIN (1,6) #13 2213 2212 2211 2210
wire n476; //IPIN (1,6) #14 452
wire n477; //IPIN (1,6) #15 453
wire n478; //OPIN (1,6) #16 2217 2216 2215 2214
wire n479; //IPIN (1,6) #17 455
wire n480; //IPIN (1,6) #18 456
wire n481; //OPIN (1,6) #19 2221 2220 2219 2218
wire n482; //IPIN (1,6) #20 458
wire n483; //IPIN (1,6) #21 459
wire n484; //OPIN (1,6) #22 2225 2224 2223 2222
wire n485; //IPIN (1,6) #23 461
wire n510; //IPIN (2,0) #0 486
wire n511; //OPIN (2,0) #1 1733 1732 1731 1730
wire n512; //IPIN (2,0) #2 488
wire n513; //IPIN (2,0) #3 489
wire n514; //OPIN (2,0) #4 1737 1736 1735 1734
wire n515; //IPIN (2,0) #5 491
wire n516; //IPIN (2,0) #6 492
wire n517; //OPIN (2,0) #7 1741 1740 1739 1738
wire n518; //IPIN (2,0) #8 494
wire n519; //IPIN (2,0) #9 495
wire n520; //OPIN (2,0) #10 1745 1744 1743 1742
wire n521; //IPIN (2,0) #11 497
wire n522; //IPIN (2,0) #12 498
wire n523; //OPIN (2,0) #13 1749 1748 1747 1746
wire n524; //IPIN (2,0) #14 500
wire n525; //IPIN (2,0) #15 501
wire n526; //OPIN (2,0) #16 1733 1732 1731 1730
wire n527; //IPIN (2,0) #17 503
wire n528; //IPIN (2,0) #18 504
wire n529; //OPIN (2,0) #19 1737 1736 1735 1734
wire n530; //IPIN (2,0) #20 506
wire n531; //IPIN (2,0) #21 507
wire n532; //OPIN (2,0) #22 1741 1740 1739 1738
wire n533; //IPIN (2,0) #23 509
wire n549; //IPIN (2,1) #0 534
wire n550; //IPIN (2,1) #1 535
wire n551; //IPIN (2,1) #2 536
wire n552; //IPIN (2,1) #3 537
wire n553; //IPIN (2,1) #4 538
wire n554; //IPIN (2,1) #5 539
wire n555; //IPIN (2,1) #6 540
wire n556; //IPIN (2,1) #7 541
wire n557; //IPIN (2,1) #8 542
wire n558; //IPIN (2,1) #9 543
wire n559; //IPIN (2,1) #10 544
wire n560; //IPIN (2,1) #11 545
wire n561; //OPIN (2,1) #12 1833 1832 1831 1830
wire n562; //OPIN (2,1) #13 2513 2512 2511 2510
wire n563; //IPIN (2,1) #14 548
wire n579; //IPIN (2,2) #0 564
wire n580; //IPIN (2,2) #1 565
wire n581; //IPIN (2,2) #2 566
wire n582; //IPIN (2,2) #3 567
wire n583; //IPIN (2,2) #4 568
wire n584; //IPIN (2,2) #5 569
wire n585; //IPIN (2,2) #6 570
wire n586; //IPIN (2,2) #7 571
wire n587; //IPIN (2,2) #8 572
wire n588; //IPIN (2,2) #9 573
wire n589; //IPIN (2,2) #10 574
wire n590; //IPIN (2,2) #11 575
wire n591; //OPIN (2,2) #12 1933 1932 1931 1930
wire n592; //OPIN (2,2) #13 2533 2532 2531 2530
wire n593; //IPIN (2,2) #14 578
wire n609; //IPIN (2,3) #0 594
wire n610; //IPIN (2,3) #1 595
wire n611; //IPIN (2,3) #2 596
wire n612; //IPIN (2,3) #3 597
wire n613; //IPIN (2,3) #4 598
wire n614; //IPIN (2,3) #5 599
wire n615; //IPIN (2,3) #6 600
wire n616; //IPIN (2,3) #7 601
wire n617; //IPIN (2,3) #8 602
wire n618; //IPIN (2,3) #9 603
wire n619; //IPIN (2,3) #10 604
wire n620; //IPIN (2,3) #11 605
wire n621; //OPIN (2,3) #12 2033 2032 2031 2030
wire n622; //OPIN (2,3) #13 2553 2552 2551 2550
wire n623; //IPIN (2,3) #14 608
wire n639; //IPIN (2,4) #0 624
wire n640; //IPIN (2,4) #1 625
wire n641; //IPIN (2,4) #2 626
wire n642; //IPIN (2,4) #3 627
wire n643; //IPIN (2,4) #4 628
wire n644; //IPIN (2,4) #5 629
wire n645; //IPIN (2,4) #6 630
wire n646; //IPIN (2,4) #7 631
wire n647; //IPIN (2,4) #8 632
wire n648; //IPIN (2,4) #9 633
wire n649; //IPIN (2,4) #10 634
wire n650; //IPIN (2,4) #11 635
wire n651; //OPIN (2,4) #12 2133 2132 2131 2130
wire n652; //OPIN (2,4) #13 2573 2572 2571 2570
wire n653; //IPIN (2,4) #14 638
wire n669; //IPIN (2,5) #0 654
wire n670; //IPIN (2,5) #1 655
wire n671; //IPIN (2,5) #2 656
wire n672; //IPIN (2,5) #3 657
wire n673; //IPIN (2,5) #4 658
wire n674; //IPIN (2,5) #5 659
wire n675; //IPIN (2,5) #6 660
wire n676; //IPIN (2,5) #7 661
wire n677; //IPIN (2,5) #8 662
wire n678; //IPIN (2,5) #9 663
wire n679; //IPIN (2,5) #10 664
wire n680; //IPIN (2,5) #11 665
wire n681; //OPIN (2,5) #12 2233 2232 2231 2230
wire n682; //OPIN (2,5) #13 2593 2592 2591 2590
wire n683; //IPIN (2,5) #14 668
wire n708; //IPIN (2,6) #0 684
wire n709; //OPIN (2,6) #1 2237 2236 2235 2234
wire n710; //IPIN (2,6) #2 686
wire n711; //IPIN (2,6) #3 687
wire n712; //OPIN (2,6) #4 2241 2240 2239 2238
wire n713; //IPIN (2,6) #5 689
wire n714; //IPIN (2,6) #6 690
wire n715; //OPIN (2,6) #7 2245 2244 2243 2242
wire n716; //IPIN (2,6) #8 692
wire n717; //IPIN (2,6) #9 693
wire n718; //OPIN (2,6) #10 2249 2248 2247 2246
wire n719; //IPIN (2,6) #11 695
wire n720; //IPIN (2,6) #12 696
wire n721; //OPIN (2,6) #13 2233 2232 2231 2230
wire n722; //IPIN (2,6) #14 698
wire n723; //IPIN (2,6) #15 699
wire n724; //OPIN (2,6) #16 2237 2236 2235 2234
wire n725; //IPIN (2,6) #17 701
wire n726; //IPIN (2,6) #18 702
wire n727; //OPIN (2,6) #19 2241 2240 2239 2238
wire n728; //IPIN (2,6) #20 704
wire n729; //IPIN (2,6) #21 705
wire n730; //OPIN (2,6) #22 2245 2244 2243 2242
wire n731; //IPIN (2,6) #23 707
wire n756; //IPIN (3,0) #0 732
wire n757; //OPIN (3,0) #1 1753 1752 1751 1750
wire n758; //IPIN (3,0) #2 734
wire n759; //IPIN (3,0) #3 735
wire n760; //OPIN (3,0) #4 1757 1756 1755 1754
wire n761; //IPIN (3,0) #5 737
wire n762; //IPIN (3,0) #6 738
wire n763; //OPIN (3,0) #7 1761 1760 1759 1758
wire n764; //IPIN (3,0) #8 740
wire n765; //IPIN (3,0) #9 741
wire n766; //OPIN (3,0) #10 1765 1764 1763 1762
wire n767; //IPIN (3,0) #11 743
wire n768; //IPIN (3,0) #12 744
wire n769; //OPIN (3,0) #13 1769 1768 1767 1766
wire n770; //IPIN (3,0) #14 746
wire n771; //IPIN (3,0) #15 747
wire n772; //OPIN (3,0) #16 1753 1752 1751 1750
wire n773; //IPIN (3,0) #17 749
wire n774; //IPIN (3,0) #18 750
wire n775; //OPIN (3,0) #19 1757 1756 1755 1754
wire n776; //IPIN (3,0) #20 752
wire n777; //IPIN (3,0) #21 753
wire n778; //OPIN (3,0) #22 1761 1760 1759 1758
wire n779; //IPIN (3,0) #23 755
wire n795; //IPIN (3,1) #0 780
wire n796; //IPIN (3,1) #1 781
wire n797; //IPIN (3,1) #2 782
wire n798; //IPIN (3,1) #3 783
wire n799; //IPIN (3,1) #4 784
wire n800; //IPIN (3,1) #5 785
wire n801; //IPIN (3,1) #6 786
wire n802; //IPIN (3,1) #7 787
wire n803; //IPIN (3,1) #8 788
wire n804; //IPIN (3,1) #9 789
wire n805; //IPIN (3,1) #10 790
wire n806; //IPIN (3,1) #11 791
wire n807; //OPIN (3,1) #12 1853 1852 1851 1850
wire n808; //OPIN (3,1) #13 2613 2612 2611 2610
wire n809; //IPIN (3,1) #14 794
wire n825; //IPIN (3,2) #0 810
wire n826; //IPIN (3,2) #1 811
wire n827; //IPIN (3,2) #2 812
wire n828; //IPIN (3,2) #3 813
wire n829; //IPIN (3,2) #4 814
wire n830; //IPIN (3,2) #5 815
wire n831; //IPIN (3,2) #6 816
wire n832; //IPIN (3,2) #7 817
wire n833; //IPIN (3,2) #8 818
wire n834; //IPIN (3,2) #9 819
wire n835; //IPIN (3,2) #10 820
wire n836; //IPIN (3,2) #11 821
wire n837; //OPIN (3,2) #12 1953 1952 1951 1950
wire n838; //OPIN (3,2) #13 2633 2632 2631 2630
wire n839; //IPIN (3,2) #14 824
wire n855; //IPIN (3,3) #0 840
wire n856; //IPIN (3,3) #1 841
wire n857; //IPIN (3,3) #2 842
wire n858; //IPIN (3,3) #3 843
wire n859; //IPIN (3,3) #4 844
wire n860; //IPIN (3,3) #5 845
wire n861; //IPIN (3,3) #6 846
wire n862; //IPIN (3,3) #7 847
wire n863; //IPIN (3,3) #8 848
wire n864; //IPIN (3,3) #9 849
wire n865; //IPIN (3,3) #10 850
wire n866; //IPIN (3,3) #11 851
wire n867; //OPIN (3,3) #12 2053 2052 2051 2050
wire n868; //OPIN (3,3) #13 2653 2652 2651 2650
wire n869; //IPIN (3,3) #14 854
wire n885; //IPIN (3,4) #0 870
wire n886; //IPIN (3,4) #1 871
wire n887; //IPIN (3,4) #2 872
wire n888; //IPIN (3,4) #3 873
wire n889; //IPIN (3,4) #4 874
wire n890; //IPIN (3,4) #5 875
wire n891; //IPIN (3,4) #6 876
wire n892; //IPIN (3,4) #7 877
wire n893; //IPIN (3,4) #8 878
wire n894; //IPIN (3,4) #9 879
wire n895; //IPIN (3,4) #10 880
wire n896; //IPIN (3,4) #11 881
wire n897; //OPIN (3,4) #12 2153 2152 2151 2150
wire n898; //OPIN (3,4) #13 2673 2672 2671 2670
wire n899; //IPIN (3,4) #14 884
wire n915; //IPIN (3,5) #0 900
wire n916; //IPIN (3,5) #1 901
wire n917; //IPIN (3,5) #2 902
wire n918; //IPIN (3,5) #3 903
wire n919; //IPIN (3,5) #4 904
wire n920; //IPIN (3,5) #5 905
wire n921; //IPIN (3,5) #6 906
wire n922; //IPIN (3,5) #7 907
wire n923; //IPIN (3,5) #8 908
wire n924; //IPIN (3,5) #9 909
wire n925; //IPIN (3,5) #10 910
wire n926; //IPIN (3,5) #11 911
wire n927; //OPIN (3,5) #12 2253 2252 2251 2250
wire n928; //OPIN (3,5) #13 2693 2692 2691 2690
wire n929; //IPIN (3,5) #14 914
wire n954; //IPIN (3,6) #0 930
wire n955; //OPIN (3,6) #1 2257 2256 2255 2254
wire n956; //IPIN (3,6) #2 932
wire n957; //IPIN (3,6) #3 933
wire n958; //OPIN (3,6) #4 2261 2260 2259 2258
wire n959; //IPIN (3,6) #5 935
wire n960; //IPIN (3,6) #6 936
wire n961; //OPIN (3,6) #7 2265 2264 2263 2262
wire n962; //IPIN (3,6) #8 938
wire n963; //IPIN (3,6) #9 939
wire n964; //OPIN (3,6) #10 2269 2268 2267 2266
wire n965; //IPIN (3,6) #11 941
wire n966; //IPIN (3,6) #12 942
wire n967; //OPIN (3,6) #13 2253 2252 2251 2250
wire n968; //IPIN (3,6) #14 944
wire n969; //IPIN (3,6) #15 945
wire n970; //OPIN (3,6) #16 2257 2256 2255 2254
wire n971; //IPIN (3,6) #17 947
wire n972; //IPIN (3,6) #18 948
wire n973; //OPIN (3,6) #19 2261 2260 2259 2258
wire n974; //IPIN (3,6) #20 950
wire n975; //IPIN (3,6) #21 951
wire n976; //OPIN (3,6) #22 2265 2264 2263 2262
wire n977; //IPIN (3,6) #23 953
wire n1002; //IPIN (4,0) #0 978
wire n1003; //OPIN (4,0) #1 1773 1772 1771 1770
wire n1004; //IPIN (4,0) #2 980
wire n1005; //IPIN (4,0) #3 981
wire n1006; //OPIN (4,0) #4 1777 1776 1775 1774
wire n1007; //IPIN (4,0) #5 983
wire n1008; //IPIN (4,0) #6 984
wire n1009; //OPIN (4,0) #7 1781 1780 1779 1778
wire n1010; //IPIN (4,0) #8 986
wire n1011; //IPIN (4,0) #9 987
wire n1012; //OPIN (4,0) #10 1785 1784 1783 1782
wire n1013; //IPIN (4,0) #11 989
wire n1014; //IPIN (4,0) #12 990
wire n1015; //OPIN (4,0) #13 1789 1788 1787 1786
wire n1016; //IPIN (4,0) #14 992
wire n1017; //IPIN (4,0) #15 993
wire n1018; //OPIN (4,0) #16 1773 1772 1771 1770
wire n1019; //IPIN (4,0) #17 995
wire n1020; //IPIN (4,0) #18 996
wire n1021; //OPIN (4,0) #19 1777 1776 1775 1774
wire n1022; //IPIN (4,0) #20 998
wire n1023; //IPIN (4,0) #21 999
wire n1024; //OPIN (4,0) #22 1781 1780 1779 1778
wire n1025; //IPIN (4,0) #23 1001
wire n1041; //IPIN (4,1) #0 1026
wire n1042; //IPIN (4,1) #1 1027
wire n1043; //IPIN (4,1) #2 1028
wire n1044; //IPIN (4,1) #3 1029
wire n1045; //IPIN (4,1) #4 1030
wire n1046; //IPIN (4,1) #5 1031
wire n1047; //IPIN (4,1) #6 1032
wire n1048; //IPIN (4,1) #7 1033
wire n1049; //IPIN (4,1) #8 1034
wire n1050; //IPIN (4,1) #9 1035
wire n1051; //IPIN (4,1) #10 1036
wire n1052; //IPIN (4,1) #11 1037
wire n1053; //OPIN (4,1) #12 1873 1872 1871 1870
wire n1054; //OPIN (4,1) #13 2713 2712 2711 2710
wire n1055; //IPIN (4,1) #14 1040
wire n1071; //IPIN (4,2) #0 1056
wire n1072; //IPIN (4,2) #1 1057
wire n1073; //IPIN (4,2) #2 1058
wire n1074; //IPIN (4,2) #3 1059
wire n1075; //IPIN (4,2) #4 1060
wire n1076; //IPIN (4,2) #5 1061
wire n1077; //IPIN (4,2) #6 1062
wire n1078; //IPIN (4,2) #7 1063
wire n1079; //IPIN (4,2) #8 1064
wire n1080; //IPIN (4,2) #9 1065
wire n1081; //IPIN (4,2) #10 1066
wire n1082; //IPIN (4,2) #11 1067
wire n1083; //OPIN (4,2) #12 1973 1972 1971 1970
wire n1084; //OPIN (4,2) #13 2733 2732 2731 2730
wire n1085; //IPIN (4,2) #14 1070
wire n1101; //IPIN (4,3) #0 1086
wire n1102; //IPIN (4,3) #1 1087
wire n1103; //IPIN (4,3) #2 1088
wire n1104; //IPIN (4,3) #3 1089
wire n1105; //IPIN (4,3) #4 1090
wire n1106; //IPIN (4,3) #5 1091
wire n1107; //IPIN (4,3) #6 1092
wire n1108; //IPIN (4,3) #7 1093
wire n1109; //IPIN (4,3) #8 1094
wire n1110; //IPIN (4,3) #9 1095
wire n1111; //IPIN (4,3) #10 1096
wire n1112; //IPIN (4,3) #11 1097
wire n1113; //OPIN (4,3) #12 2073 2072 2071 2070
wire n1114; //OPIN (4,3) #13 2753 2752 2751 2750
wire n1115; //IPIN (4,3) #14 1100
wire n1131; //IPIN (4,4) #0 1116
wire n1132; //IPIN (4,4) #1 1117
wire n1133; //IPIN (4,4) #2 1118
wire n1134; //IPIN (4,4) #3 1119
wire n1135; //IPIN (4,4) #4 1120
wire n1136; //IPIN (4,4) #5 1121
wire n1137; //IPIN (4,4) #6 1122
wire n1138; //IPIN (4,4) #7 1123
wire n1139; //IPIN (4,4) #8 1124
wire n1140; //IPIN (4,4) #9 1125
wire n1141; //IPIN (4,4) #10 1126
wire n1142; //IPIN (4,4) #11 1127
wire n1143; //OPIN (4,4) #12 2173 2172 2171 2170
wire n1144; //OPIN (4,4) #13 2773 2772 2771 2770
wire n1145; //IPIN (4,4) #14 1130
wire n1161; //IPIN (4,5) #0 1146
wire n1162; //IPIN (4,5) #1 1147
wire n1163; //IPIN (4,5) #2 1148
wire n1164; //IPIN (4,5) #3 1149
wire n1165; //IPIN (4,5) #4 1150
wire n1166; //IPIN (4,5) #5 1151
wire n1167; //IPIN (4,5) #6 1152
wire n1168; //IPIN (4,5) #7 1153
wire n1169; //IPIN (4,5) #8 1154
wire n1170; //IPIN (4,5) #9 1155
wire n1171; //IPIN (4,5) #10 1156
wire n1172; //IPIN (4,5) #11 1157
wire n1173; //OPIN (4,5) #12 2273 2272 2271 2270
wire n1174; //OPIN (4,5) #13 2793 2792 2791 2790
wire n1175; //IPIN (4,5) #14 1160
wire n1200; //IPIN (4,6) #0 1176
wire n1201; //OPIN (4,6) #1 2277 2276 2275 2274
wire n1202; //IPIN (4,6) #2 1178
wire n1203; //IPIN (4,6) #3 1179
wire n1204; //OPIN (4,6) #4 2281 2280 2279 2278
wire n1205; //IPIN (4,6) #5 1181
wire n1206; //IPIN (4,6) #6 1182
wire n1207; //OPIN (4,6) #7 2285 2284 2283 2282
wire n1208; //IPIN (4,6) #8 1184
wire n1209; //IPIN (4,6) #9 1185
wire n1210; //OPIN (4,6) #10 2289 2288 2287 2286
wire n1211; //IPIN (4,6) #11 1187
wire n1212; //IPIN (4,6) #12 1188
wire n1213; //OPIN (4,6) #13 2273 2272 2271 2270
wire n1214; //IPIN (4,6) #14 1190
wire n1215; //IPIN (4,6) #15 1191
wire n1216; //OPIN (4,6) #16 2277 2276 2275 2274
wire n1217; //IPIN (4,6) #17 1193
wire n1218; //IPIN (4,6) #18 1194
wire n1219; //OPIN (4,6) #19 2281 2280 2279 2278
wire n1220; //IPIN (4,6) #20 1196
wire n1221; //IPIN (4,6) #21 1197
wire n1222; //OPIN (4,6) #22 2285 2284 2283 2282
wire n1223; //IPIN (4,6) #23 1199
wire n1248; //IPIN (5,0) #0 1224
wire n1249; //OPIN (5,0) #1 1793 1792 1791 1790
wire n1250; //IPIN (5,0) #2 1226
wire n1251; //IPIN (5,0) #3 1227
wire n1252; //OPIN (5,0) #4 1797 1796 1795 1794
wire n1253; //IPIN (5,0) #5 1229
wire n1254; //IPIN (5,0) #6 1230
wire n1255; //OPIN (5,0) #7 1801 1800 1799 1798
wire n1256; //IPIN (5,0) #8 1232
wire n1257; //IPIN (5,0) #9 1233
wire n1258; //OPIN (5,0) #10 1805 1804 1803 1802
wire n1259; //IPIN (5,0) #11 1235
wire n1260; //IPIN (5,0) #12 1236
wire n1261; //OPIN (5,0) #13 1809 1808 1807 1806
wire n1262; //IPIN (5,0) #14 1238
wire n1263; //IPIN (5,0) #15 1239
wire n1264; //OPIN (5,0) #16 1793 1792 1791 1790
wire n1265; //IPIN (5,0) #17 1241
wire n1266; //IPIN (5,0) #18 1242
wire n1267; //OPIN (5,0) #19 1797 1796 1795 1794
wire n1268; //IPIN (5,0) #20 1244
wire n1269; //IPIN (5,0) #21 1245
wire n1270; //OPIN (5,0) #22 1801 1800 1799 1798
wire n1271; //IPIN (5,0) #23 1247
wire n1287; //IPIN (5,1) #0 1272
wire n1288; //IPIN (5,1) #1 1273
wire n1289; //IPIN (5,1) #2 1274
wire n1290; //IPIN (5,1) #3 1275
wire n1291; //IPIN (5,1) #4 1276
wire n1292; //IPIN (5,1) #5 1277
wire n1293; //IPIN (5,1) #6 1278
wire n1294; //IPIN (5,1) #7 1279
wire n1295; //IPIN (5,1) #8 1280
wire n1296; //IPIN (5,1) #9 1281
wire n1297; //IPIN (5,1) #10 1282
wire n1298; //IPIN (5,1) #11 1283
wire n1299; //OPIN (5,1) #12 1893 1892 1891 1890
wire n1300; //OPIN (5,1) #13 2813 2812 2811 2810
wire n1301; //IPIN (5,1) #14 1286
wire n1317; //IPIN (5,2) #0 1302
wire n1318; //IPIN (5,2) #1 1303
wire n1319; //IPIN (5,2) #2 1304
wire n1320; //IPIN (5,2) #3 1305
wire n1321; //IPIN (5,2) #4 1306
wire n1322; //IPIN (5,2) #5 1307
wire n1323; //IPIN (5,2) #6 1308
wire n1324; //IPIN (5,2) #7 1309
wire n1325; //IPIN (5,2) #8 1310
wire n1326; //IPIN (5,2) #9 1311
wire n1327; //IPIN (5,2) #10 1312
wire n1328; //IPIN (5,2) #11 1313
wire n1329; //OPIN (5,2) #12 1993 1992 1991 1990
wire n1330; //OPIN (5,2) #13 2833 2832 2831 2830
wire n1331; //IPIN (5,2) #14 1316
wire n1347; //IPIN (5,3) #0 1332
wire n1348; //IPIN (5,3) #1 1333
wire n1349; //IPIN (5,3) #2 1334
wire n1350; //IPIN (5,3) #3 1335
wire n1351; //IPIN (5,3) #4 1336
wire n1352; //IPIN (5,3) #5 1337
wire n1353; //IPIN (5,3) #6 1338
wire n1354; //IPIN (5,3) #7 1339
wire n1355; //IPIN (5,3) #8 1340
wire n1356; //IPIN (5,3) #9 1341
wire n1357; //IPIN (5,3) #10 1342
wire n1358; //IPIN (5,3) #11 1343
wire n1359; //OPIN (5,3) #12 2093 2092 2091 2090
wire n1360; //OPIN (5,3) #13 2853 2852 2851 2850
wire n1361; //IPIN (5,3) #14 1346
wire n1377; //IPIN (5,4) #0 1362
wire n1378; //IPIN (5,4) #1 1363
wire n1379; //IPIN (5,4) #2 1364
wire n1380; //IPIN (5,4) #3 1365
wire n1381; //IPIN (5,4) #4 1366
wire n1382; //IPIN (5,4) #5 1367
wire n1383; //IPIN (5,4) #6 1368
wire n1384; //IPIN (5,4) #7 1369
wire n1385; //IPIN (5,4) #8 1370
wire n1386; //IPIN (5,4) #9 1371
wire n1387; //IPIN (5,4) #10 1372
wire n1388; //IPIN (5,4) #11 1373
wire n1389; //OPIN (5,4) #12 2193 2192 2191 2190
wire n1390; //OPIN (5,4) #13 2873 2872 2871 2870
wire n1391; //IPIN (5,4) #14 1376
wire n1407; //IPIN (5,5) #0 1392
wire n1408; //IPIN (5,5) #1 1393
wire n1409; //IPIN (5,5) #2 1394
wire n1410; //IPIN (5,5) #3 1395
wire n1411; //IPIN (5,5) #4 1396
wire n1412; //IPIN (5,5) #5 1397
wire n1413; //IPIN (5,5) #6 1398
wire n1414; //IPIN (5,5) #7 1399
wire n1415; //IPIN (5,5) #8 1400
wire n1416; //IPIN (5,5) #9 1401
wire n1417; //IPIN (5,5) #10 1402
wire n1418; //IPIN (5,5) #11 1403
wire n1419; //OPIN (5,5) #12 2293 2292 2291 2290
wire n1420; //OPIN (5,5) #13 2893 2892 2891 2890
wire n1421; //IPIN (5,5) #14 1406
wire n1446; //IPIN (5,6) #0 1422
wire n1447; //OPIN (5,6) #1 2297 2296 2295 2294
wire n1448; //IPIN (5,6) #2 1424
wire n1449; //IPIN (5,6) #3 1425
wire n1450; //OPIN (5,6) #4 2301 2300 2299 2298
wire n1451; //IPIN (5,6) #5 1427
wire n1452; //IPIN (5,6) #6 1428
wire n1453; //OPIN (5,6) #7 2305 2304 2303 2302
wire n1454; //IPIN (5,6) #8 1430
wire n1455; //IPIN (5,6) #9 1431
wire n1456; //OPIN (5,6) #10 2309 2308 2307 2306
wire n1457; //IPIN (5,6) #11 1433
wire n1458; //IPIN (5,6) #12 1434
wire n1459; //OPIN (5,6) #13 2293 2292 2291 2290
wire n1460; //IPIN (5,6) #14 1436
wire n1461; //IPIN (5,6) #15 1437
wire n1462; //OPIN (5,6) #16 2297 2296 2295 2294
wire n1463; //IPIN (5,6) #17 1439
wire n1464; //IPIN (5,6) #18 1440
wire n1465; //OPIN (5,6) #19 2301 2300 2299 2298
wire n1466; //IPIN (5,6) #20 1442
wire n1467; //IPIN (5,6) #21 1443
wire n1468; //OPIN (5,6) #22 2305 2304 2303 2302
wire n1469; //IPIN (5,6) #23 1445
wire n1494; //IPIN (6,1) #0 1470
wire n1495; //OPIN (6,1) #1 2817 2816 2815 2814
wire n1496; //IPIN (6,1) #2 1472
wire n1497; //IPIN (6,1) #3 1473
wire n1498; //OPIN (6,1) #4 2821 2820 2819 2818
wire n1499; //IPIN (6,1) #5 1475
wire n1500; //IPIN (6,1) #6 1476
wire n1501; //OPIN (6,1) #7 2825 2824 2823 2822
wire n1502; //IPIN (6,1) #8 1478
wire n1503; //IPIN (6,1) #9 1479
wire n1504; //OPIN (6,1) #10 2829 2828 2827 2826
wire n1505; //IPIN (6,1) #11 1481
wire n1506; //IPIN (6,1) #12 1482
wire n1507; //OPIN (6,1) #13 2813 2812 2811 2810
wire n1508; //IPIN (6,1) #14 1484
wire n1509; //IPIN (6,1) #15 1485
wire n1510; //OPIN (6,1) #16 2817 2816 2815 2814
wire n1511; //IPIN (6,1) #17 1487
wire n1512; //IPIN (6,1) #18 1488
wire n1513; //OPIN (6,1) #19 2821 2820 2819 2818
wire n1514; //IPIN (6,1) #20 1490
wire n1515; //IPIN (6,1) #21 1491
wire n1516; //OPIN (6,1) #22 2825 2824 2823 2822
wire n1517; //IPIN (6,1) #23 1493
wire n1542; //IPIN (6,2) #0 1518
wire n1543; //OPIN (6,2) #1 2837 2836 2835 2834
wire n1544; //IPIN (6,2) #2 1520
wire n1545; //IPIN (6,2) #3 1521
wire n1546; //OPIN (6,2) #4 2841 2840 2839 2838
wire n1547; //IPIN (6,2) #5 1523
wire n1548; //IPIN (6,2) #6 1524
wire n1549; //OPIN (6,2) #7 2845 2844 2843 2842
wire n1550; //IPIN (6,2) #8 1526
wire n1551; //IPIN (6,2) #9 1527
wire n1552; //OPIN (6,2) #10 2849 2848 2847 2846
wire n1553; //IPIN (6,2) #11 1529
wire n1554; //IPIN (6,2) #12 1530
wire n1555; //OPIN (6,2) #13 2833 2832 2831 2830
wire n1556; //IPIN (6,2) #14 1532
wire n1557; //IPIN (6,2) #15 1533
wire n1558; //OPIN (6,2) #16 2837 2836 2835 2834
wire n1559; //IPIN (6,2) #17 1535
wire n1560; //IPIN (6,2) #18 1536
wire n1561; //OPIN (6,2) #19 2841 2840 2839 2838
wire n1562; //IPIN (6,2) #20 1538
wire n1563; //IPIN (6,2) #21 1539
wire n1564; //OPIN (6,2) #22 2845 2844 2843 2842
wire n1565; //IPIN (6,2) #23 1541
wire n1590; //IPIN (6,3) #0 1566
wire n1591; //OPIN (6,3) #1 2857 2856 2855 2854
wire n1592; //IPIN (6,3) #2 1568
wire n1593; //IPIN (6,3) #3 1569
wire n1594; //OPIN (6,3) #4 2861 2860 2859 2858
wire n1595; //IPIN (6,3) #5 1571
wire n1596; //IPIN (6,3) #6 1572
wire n1597; //OPIN (6,3) #7 2865 2864 2863 2862
wire n1598; //IPIN (6,3) #8 1574
wire n1599; //IPIN (6,3) #9 1575
wire n1600; //OPIN (6,3) #10 2869 2868 2867 2866
wire n1601; //IPIN (6,3) #11 1577
wire n1602; //IPIN (6,3) #12 1578
wire n1603; //OPIN (6,3) #13 2853 2852 2851 2850
wire n1604; //IPIN (6,3) #14 1580
wire n1605; //IPIN (6,3) #15 1581
wire n1606; //OPIN (6,3) #16 2857 2856 2855 2854
wire n1607; //IPIN (6,3) #17 1583
wire n1608; //IPIN (6,3) #18 1584
wire n1609; //OPIN (6,3) #19 2861 2860 2859 2858
wire n1610; //IPIN (6,3) #20 1586
wire n1611; //IPIN (6,3) #21 1587
wire n1612; //OPIN (6,3) #22 2865 2864 2863 2862
wire n1613; //IPIN (6,3) #23 1589
wire n1638; //IPIN (6,4) #0 1614
wire n1639; //OPIN (6,4) #1 2877 2876 2875 2874
wire n1640; //IPIN (6,4) #2 1616
wire n1641; //IPIN (6,4) #3 1617
wire n1642; //OPIN (6,4) #4 2881 2880 2879 2878
wire n1643; //IPIN (6,4) #5 1619
wire n1644; //IPIN (6,4) #6 1620
wire n1645; //OPIN (6,4) #7 2885 2884 2883 2882
wire n1646; //IPIN (6,4) #8 1622
wire n1647; //IPIN (6,4) #9 1623
wire n1648; //OPIN (6,4) #10 2889 2888 2887 2886
wire n1649; //IPIN (6,4) #11 1625
wire n1650; //IPIN (6,4) #12 1626
wire n1651; //OPIN (6,4) #13 2873 2872 2871 2870
wire n1652; //IPIN (6,4) #14 1628
wire n1653; //IPIN (6,4) #15 1629
wire n1654; //OPIN (6,4) #16 2877 2876 2875 2874
wire n1655; //IPIN (6,4) #17 1631
wire n1656; //IPIN (6,4) #18 1632
wire n1657; //OPIN (6,4) #19 2881 2880 2879 2878
wire n1658; //IPIN (6,4) #20 1634
wire n1659; //IPIN (6,4) #21 1635
wire n1660; //OPIN (6,4) #22 2885 2884 2883 2882
wire n1661; //IPIN (6,4) #23 1637
wire n1686; //IPIN (6,5) #0 1662
wire n1687; //OPIN (6,5) #1 2897 2896 2895 2894
wire n1688; //IPIN (6,5) #2 1664
wire n1689; //IPIN (6,5) #3 1665
wire n1690; //OPIN (6,5) #4 2901 2900 2899 2898
wire n1691; //IPIN (6,5) #5 1667
wire n1692; //IPIN (6,5) #6 1668
wire n1693; //OPIN (6,5) #7 2905 2904 2903 2902
wire n1694; //IPIN (6,5) #8 1670
wire n1695; //IPIN (6,5) #9 1671
wire n1696; //OPIN (6,5) #10 2909 2908 2907 2906
wire n1697; //IPIN (6,5) #11 1673
wire n1698; //IPIN (6,5) #12 1674
wire n1699; //OPIN (6,5) #13 2893 2892 2891 2890
wire n1700; //IPIN (6,5) #14 1676
wire n1701; //IPIN (6,5) #15 1677
wire n1702; //OPIN (6,5) #16 2897 2896 2895 2894
wire n1703; //IPIN (6,5) #17 1679
wire n1704; //IPIN (6,5) #18 1680
wire n1705; //OPIN (6,5) #19 2901 2900 2899 2898
wire n1706; //IPIN (6,5) #20 1682
wire n1707; //IPIN (6,5) #21 1683
wire n1708; //OPIN (6,5) #22 2905 2904 2903 2902
wire n1709; //IPIN (6,5) #23 1685
wire n1710; //CHANX (1,0) #0 1730 2414 305 267 264
wire n1711; //CHANX (1,0) #1 2328 305 267 264
wire n1712; //CHANX (1,0) #2 1732 2420 273 270
wire n1713; //CHANX (1,0) #3 2310 273 270
wire n1714; //CHANX (1,0) #4 1734 2426 309 276
wire n1715; //CHANX (1,0) #5 2312 309 276
wire n1716; //CHANX (1,0) #6 1736 2410 282 279
wire n1717; //CHANX (1,0) #7 2314 282 279
wire n1718; //CHANX (1,0) #8 1738 2412 313 285
wire n1719; //CHANX (1,0) #9 2316 313 285
wire n1720; //CHANX (1,0) #10 1740 2416 305 267 264
wire n1721; //CHANX (1,0) #11 2318 305 267 264
wire n1722; //CHANX (1,0) #12 1742 2418 273 270
wire n1723; //CHANX (1,0) #13 2320 273 270
wire n1724; //CHANX (1,0) #14 1744 2422 309 276
wire n1725; //CHANX (1,0) #15 2322 309 276
wire n1726; //CHANX (1,0) #16 1746 2424 282 279
wire n1727; //CHANX (1,0) #17 2324 282 279
wire n1728; //CHANX (1,0) #18 1748 2428 313 285
wire n1729; //CHANX (1,0) #19 2326 313 285
wire n1730; //CHANX (2,0) #0 1750 2514 551 513 510
wire n1731; //CHANX (2,0) #1 1711 2414 551 513 510
wire n1732; //CHANX (2,0) #2 1752 2520 519 516
wire n1733; //CHANX (2,0) #3 1713 2420 519 516
wire n1734; //CHANX (2,0) #4 1754 2526 555 522
wire n1735; //CHANX (2,0) #5 1715 2426 555 522
wire n1736; //CHANX (2,0) #6 1756 2510 528 525
wire n1737; //CHANX (2,0) #7 1717 2410 528 525
wire n1738; //CHANX (2,0) #8 1758 2512 559 531
wire n1739; //CHANX (2,0) #9 1719 2412 559 531
wire n1740; //CHANX (2,0) #10 1760 2516 551 513 510
wire n1741; //CHANX (2,0) #11 1721 2416 551 513 510
wire n1742; //CHANX (2,0) #12 1762 2518 519 516
wire n1743; //CHANX (2,0) #13 1723 2418 519 516
wire n1744; //CHANX (2,0) #14 1764 2522 555 522
wire n1745; //CHANX (2,0) #15 1725 2422 555 522
wire n1746; //CHANX (2,0) #16 1766 2524 528 525
wire n1747; //CHANX (2,0) #17 1727 2424 528 525
wire n1748; //CHANX (2,0) #18 1768 2528 559 531
wire n1749; //CHANX (2,0) #19 1729 2428 559 531
wire n1750; //CHANX (3,0) #0 1770 2614 797 759 756
wire n1751; //CHANX (3,0) #1 1731 2514 797 759 756
wire n1752; //CHANX (3,0) #2 1772 2620 765 762
wire n1753; //CHANX (3,0) #3 1733 2520 765 762
wire n1754; //CHANX (3,0) #4 1774 2626 801 768
wire n1755; //CHANX (3,0) #5 1735 2526 801 768
wire n1756; //CHANX (3,0) #6 1776 2610 774 771
wire n1757; //CHANX (3,0) #7 1737 2510 774 771
wire n1758; //CHANX (3,0) #8 1778 2612 805 777
wire n1759; //CHANX (3,0) #9 1739 2512 805 777
wire n1760; //CHANX (3,0) #10 1780 2616 797 759 756
wire n1761; //CHANX (3,0) #11 1741 2516 797 759 756
wire n1762; //CHANX (3,0) #12 1782 2618 765 762
wire n1763; //CHANX (3,0) #13 1743 2518 765 762
wire n1764; //CHANX (3,0) #14 1784 2622 801 768
wire n1765; //CHANX (3,0) #15 1745 2522 801 768
wire n1766; //CHANX (3,0) #16 1786 2624 774 771
wire n1767; //CHANX (3,0) #17 1747 2524 774 771
wire n1768; //CHANX (3,0) #18 1788 2628 805 777
wire n1769; //CHANX (3,0) #19 1749 2528 805 777
wire n1770; //CHANX (4,0) #0 1790 2714 1043 1005 1002
wire n1771; //CHANX (4,0) #1 1751 2614 1043 1005 1002
wire n1772; //CHANX (4,0) #2 1792 2720 1011 1008
wire n1773; //CHANX (4,0) #3 1753 2620 1011 1008
wire n1774; //CHANX (4,0) #4 1794 2726 1047 1014
wire n1775; //CHANX (4,0) #5 1755 2626 1047 1014
wire n1776; //CHANX (4,0) #6 1796 2710 1020 1017
wire n1777; //CHANX (4,0) #7 1757 2610 1020 1017
wire n1778; //CHANX (4,0) #8 1798 2712 1051 1023
wire n1779; //CHANX (4,0) #9 1759 2612 1051 1023
wire n1780; //CHANX (4,0) #10 1800 2716 1043 1005 1002
wire n1781; //CHANX (4,0) #11 1761 2616 1043 1005 1002
wire n1782; //CHANX (4,0) #12 1802 2718 1011 1008
wire n1783; //CHANX (4,0) #13 1763 2618 1011 1008
wire n1784; //CHANX (4,0) #14 1804 2722 1047 1014
wire n1785; //CHANX (4,0) #15 1765 2622 1047 1014
wire n1786; //CHANX (4,0) #16 1806 2724 1020 1017
wire n1787; //CHANX (4,0) #17 1767 2624 1020 1017
wire n1788; //CHANX (4,0) #18 1808 2728 1051 1023
wire n1789; //CHANX (4,0) #19 1769 2628 1051 1023
wire n1790; //CHANX (5,0) #0 2810 1289 1251 1248
wire n1791; //CHANX (5,0) #1 1771 2714 1289 1251 1248
wire n1792; //CHANX (5,0) #2 2828 1257 1254
wire n1793; //CHANX (5,0) #3 1773 2720 1257 1254
wire n1794; //CHANX (5,0) #4 2826 1293 1260
wire n1795; //CHANX (5,0) #5 1775 2726 1293 1260
wire n1796; //CHANX (5,0) #6 2824 1266 1263
wire n1797; //CHANX (5,0) #7 1777 2710 1266 1263
wire n1798; //CHANX (5,0) #8 2822 1297 1269
wire n1799; //CHANX (5,0) #9 1779 2712 1297 1269
wire n1800; //CHANX (5,0) #10 2820 1289 1251 1248
wire n1801; //CHANX (5,0) #11 1781 2716 1289 1251 1248
wire n1802; //CHANX (5,0) #12 2818 1257 1254
wire n1803; //CHANX (5,0) #13 1783 2718 1257 1254
wire n1804; //CHANX (5,0) #14 2816 1293 1260
wire n1805; //CHANX (5,0) #15 1785 2722 1293 1260
wire n1806; //CHANX (5,0) #16 2814 1266 1263
wire n1807; //CHANX (5,0) #17 1787 2724 1266 1263
wire n1808; //CHANX (5,0) #18 2812 1297 1269
wire n1809; //CHANX (5,0) #19 1789 2728 1297 1269
wire n1810; //CHANX (1,1) #0 1830 2430 2429 335 303
wire n1811; //CHANX (1,1) #1 2330 2311 335 303
wire n1812; //CHANX (1,1) #2 1832 2448 2411 307
wire n1813; //CHANX (1,1) #3 2332 2313 307
wire n1814; //CHANX (1,1) #4 1834 2446 2413 339
wire n1815; //CHANX (1,1) #5 2334 2315 339
wire n1816; //CHANX (1,1) #6 1836 2444 2415 311
wire n1817; //CHANX (1,1) #7 2336 2317 311
wire n1818; //CHANX (1,1) #8 1838 2442 2417 343
wire n1819; //CHANX (1,1) #9 2338 2319 343
wire n1820; //CHANX (1,1) #10 1840 2440 2419 335 303
wire n1821; //CHANX (1,1) #11 2340 2321 335 303
wire n1822; //CHANX (1,1) #12 1842 2438 2421 307
wire n1823; //CHANX (1,1) #13 2342 2323 307
wire n1824; //CHANX (1,1) #14 1844 2436 2423 339
wire n1825; //CHANX (1,1) #15 2344 2325 339
wire n1826; //CHANX (1,1) #16 1846 2434 2425 311
wire n1827; //CHANX (1,1) #17 2346 2327 311
wire n1828; //CHANX (1,1) #18 1848 2432 2427 343
wire n1829; //CHANX (1,1) #19 2348 2329 343
wire n1830; //CHANX (2,1) #0 1850 2530 2529 581 549
wire n1831; //CHANX (2,1) #1 1811 2448 2427 581 549
wire n1832; //CHANX (2,1) #2 1852 2548 2511 553
wire n1833; //CHANX (2,1) #3 1813 2430 2425 553
wire n1834; //CHANX (2,1) #4 1854 2546 2513 585
wire n1835; //CHANX (2,1) #5 1815 2432 2423 585
wire n1836; //CHANX (2,1) #6 1856 2544 2515 557
wire n1837; //CHANX (2,1) #7 1817 2434 2421 557
wire n1838; //CHANX (2,1) #8 1858 2542 2517 589
wire n1839; //CHANX (2,1) #9 1819 2436 2419 589
wire n1840; //CHANX (2,1) #10 1860 2540 2519 581 549
wire n1841; //CHANX (2,1) #11 1821 2438 2417 581 549
wire n1842; //CHANX (2,1) #12 1862 2538 2521 553
wire n1843; //CHANX (2,1) #13 1823 2440 2415 553
wire n1844; //CHANX (2,1) #14 1864 2536 2523 585
wire n1845; //CHANX (2,1) #15 1825 2442 2413 585
wire n1846; //CHANX (2,1) #16 1866 2534 2525 557
wire n1847; //CHANX (2,1) #17 1827 2444 2411 557
wire n1848; //CHANX (2,1) #18 1868 2532 2527 589
wire n1849; //CHANX (2,1) #19 1829 2446 2429 589
wire n1850; //CHANX (3,1) #0 1870 2630 2629 827 795
wire n1851; //CHANX (3,1) #1 1831 2548 2527 827 795
wire n1852; //CHANX (3,1) #2 1872 2648 2611 799
wire n1853; //CHANX (3,1) #3 1833 2530 2525 799
wire n1854; //CHANX (3,1) #4 1874 2646 2613 831
wire n1855; //CHANX (3,1) #5 1835 2532 2523 831
wire n1856; //CHANX (3,1) #6 1876 2644 2615 803
wire n1857; //CHANX (3,1) #7 1837 2534 2521 803
wire n1858; //CHANX (3,1) #8 1878 2642 2617 835
wire n1859; //CHANX (3,1) #9 1839 2536 2519 835
wire n1860; //CHANX (3,1) #10 1880 2640 2619 827 795
wire n1861; //CHANX (3,1) #11 1841 2538 2517 827 795
wire n1862; //CHANX (3,1) #12 1882 2638 2621 799
wire n1863; //CHANX (3,1) #13 1843 2540 2515 799
wire n1864; //CHANX (3,1) #14 1884 2636 2623 831
wire n1865; //CHANX (3,1) #15 1845 2542 2513 831
wire n1866; //CHANX (3,1) #16 1886 2634 2625 803
wire n1867; //CHANX (3,1) #17 1847 2544 2511 803
wire n1868; //CHANX (3,1) #18 1888 2632 2627 835
wire n1869; //CHANX (3,1) #19 1849 2546 2529 835
wire n1870; //CHANX (4,1) #0 1890 2730 2729 1073 1041
wire n1871; //CHANX (4,1) #1 1851 2648 2627 1073 1041
wire n1872; //CHANX (4,1) #2 1892 2748 2711 1045
wire n1873; //CHANX (4,1) #3 1853 2630 2625 1045
wire n1874; //CHANX (4,1) #4 1894 2746 2713 1077
wire n1875; //CHANX (4,1) #5 1855 2632 2623 1077
wire n1876; //CHANX (4,1) #6 1896 2744 2715 1049
wire n1877; //CHANX (4,1) #7 1857 2634 2621 1049
wire n1878; //CHANX (4,1) #8 1898 2742 2717 1081
wire n1879; //CHANX (4,1) #9 1859 2636 2619 1081
wire n1880; //CHANX (4,1) #10 1900 2740 2719 1073 1041
wire n1881; //CHANX (4,1) #11 1861 2638 2617 1073 1041
wire n1882; //CHANX (4,1) #12 1902 2738 2721 1045
wire n1883; //CHANX (4,1) #13 1863 2640 2615 1045
wire n1884; //CHANX (4,1) #14 1904 2736 2723 1077
wire n1885; //CHANX (4,1) #15 1865 2642 2613 1077
wire n1886; //CHANX (4,1) #16 1906 2734 2725 1049
wire n1887; //CHANX (4,1) #17 1867 2644 2611 1049
wire n1888; //CHANX (4,1) #18 1908 2732 2727 1081
wire n1889; //CHANX (4,1) #19 1869 2646 2629 1081
wire n1890; //CHANX (5,1) #0 2830 2811 1319 1287
wire n1891; //CHANX (5,1) #1 1871 2748 2727 1319 1287
wire n1892; //CHANX (5,1) #2 2832 2813 1291
wire n1893; //CHANX (5,1) #3 1873 2730 2725 1291
wire n1894; //CHANX (5,1) #4 2834 2815 1323
wire n1895; //CHANX (5,1) #5 1875 2732 2723 1323
wire n1896; //CHANX (5,1) #6 2836 2817 1295
wire n1897; //CHANX (5,1) #7 1877 2734 2721 1295
wire n1898; //CHANX (5,1) #8 2838 2819 1327
wire n1899; //CHANX (5,1) #9 1879 2736 2719 1327
wire n1900; //CHANX (5,1) #10 2840 2821 1319 1287
wire n1901; //CHANX (5,1) #11 1881 2738 2717 1319 1287
wire n1902; //CHANX (5,1) #12 2842 2823 1291
wire n1903; //CHANX (5,1) #13 1883 2740 2715 1291
wire n1904; //CHANX (5,1) #14 2844 2825 1323
wire n1905; //CHANX (5,1) #15 1885 2742 2713 1323
wire n1906; //CHANX (5,1) #16 2846 2827 1295
wire n1907; //CHANX (5,1) #17 1887 2744 2711 1295
wire n1908; //CHANX (5,1) #18 2848 2829 1327
wire n1909; //CHANX (5,1) #19 1889 2746 2729 1327
wire n1910; //CHANX (1,2) #0 1930 2450 2449 365 333
wire n1911; //CHANX (1,2) #1 2350 2331 365 333
wire n1912; //CHANX (1,2) #2 1932 2468 2431 337
wire n1913; //CHANX (1,2) #3 2352 2333 337
wire n1914; //CHANX (1,2) #4 1934 2466 2433 369
wire n1915; //CHANX (1,2) #5 2354 2335 369
wire n1916; //CHANX (1,2) #6 1936 2464 2435 341
wire n1917; //CHANX (1,2) #7 2356 2337 341
wire n1918; //CHANX (1,2) #8 1938 2462 2437 373
wire n1919; //CHANX (1,2) #9 2358 2339 373
wire n1920; //CHANX (1,2) #10 1940 2460 2439 365 333
wire n1921; //CHANX (1,2) #11 2360 2341 365 333
wire n1922; //CHANX (1,2) #12 1942 2458 2441 337
wire n1923; //CHANX (1,2) #13 2362 2343 337
wire n1924; //CHANX (1,2) #14 1944 2456 2443 369
wire n1925; //CHANX (1,2) #15 2364 2345 369
wire n1926; //CHANX (1,2) #16 1946 2454 2445 341
wire n1927; //CHANX (1,2) #17 2366 2347 341
wire n1928; //CHANX (1,2) #18 1948 2452 2447 373
wire n1929; //CHANX (1,2) #19 2368 2349 373
wire n1930; //CHANX (2,2) #0 1950 2550 2549 611 579
wire n1931; //CHANX (2,2) #1 1911 2468 2447 611 579
wire n1932; //CHANX (2,2) #2 1952 2568 2531 583
wire n1933; //CHANX (2,2) #3 1913 2450 2445 583
wire n1934; //CHANX (2,2) #4 1954 2566 2533 615
wire n1935; //CHANX (2,2) #5 1915 2452 2443 615
wire n1936; //CHANX (2,2) #6 1956 2564 2535 587
wire n1937; //CHANX (2,2) #7 1917 2454 2441 587
wire n1938; //CHANX (2,2) #8 1958 2562 2537 619
wire n1939; //CHANX (2,2) #9 1919 2456 2439 619
wire n1940; //CHANX (2,2) #10 1960 2560 2539 611 579
wire n1941; //CHANX (2,2) #11 1921 2458 2437 611 579
wire n1942; //CHANX (2,2) #12 1962 2558 2541 583
wire n1943; //CHANX (2,2) #13 1923 2460 2435 583
wire n1944; //CHANX (2,2) #14 1964 2556 2543 615
wire n1945; //CHANX (2,2) #15 1925 2462 2433 615
wire n1946; //CHANX (2,2) #16 1966 2554 2545 587
wire n1947; //CHANX (2,2) #17 1927 2464 2431 587
wire n1948; //CHANX (2,2) #18 1968 2552 2547 619
wire n1949; //CHANX (2,2) #19 1929 2466 2449 619
wire n1950; //CHANX (3,2) #0 1970 2650 2649 857 825
wire n1951; //CHANX (3,2) #1 1931 2568 2547 857 825
wire n1952; //CHANX (3,2) #2 1972 2668 2631 829
wire n1953; //CHANX (3,2) #3 1933 2550 2545 829
wire n1954; //CHANX (3,2) #4 1974 2666 2633 861
wire n1955; //CHANX (3,2) #5 1935 2552 2543 861
wire n1956; //CHANX (3,2) #6 1976 2664 2635 833
wire n1957; //CHANX (3,2) #7 1937 2554 2541 833
wire n1958; //CHANX (3,2) #8 1978 2662 2637 865
wire n1959; //CHANX (3,2) #9 1939 2556 2539 865
wire n1960; //CHANX (3,2) #10 1980 2660 2639 857 825
wire n1961; //CHANX (3,2) #11 1941 2558 2537 857 825
wire n1962; //CHANX (3,2) #12 1982 2658 2641 829
wire n1963; //CHANX (3,2) #13 1943 2560 2535 829
wire n1964; //CHANX (3,2) #14 1984 2656 2643 861
wire n1965; //CHANX (3,2) #15 1945 2562 2533 861
wire n1966; //CHANX (3,2) #16 1986 2654 2645 833
wire n1967; //CHANX (3,2) #17 1947 2564 2531 833
wire n1968; //CHANX (3,2) #18 1988 2652 2647 865
wire n1969; //CHANX (3,2) #19 1949 2566 2549 865
wire n1970; //CHANX (4,2) #0 1990 2750 2749 1103 1071
wire n1971; //CHANX (4,2) #1 1951 2668 2647 1103 1071
wire n1972; //CHANX (4,2) #2 1992 2768 2731 1075
wire n1973; //CHANX (4,2) #3 1953 2650 2645 1075
wire n1974; //CHANX (4,2) #4 1994 2766 2733 1107
wire n1975; //CHANX (4,2) #5 1955 2652 2643 1107
wire n1976; //CHANX (4,2) #6 1996 2764 2735 1079
wire n1977; //CHANX (4,2) #7 1957 2654 2641 1079
wire n1978; //CHANX (4,2) #8 1998 2762 2737 1111
wire n1979; //CHANX (4,2) #9 1959 2656 2639 1111
wire n1980; //CHANX (4,2) #10 2000 2760 2739 1103 1071
wire n1981; //CHANX (4,2) #11 1961 2658 2637 1103 1071
wire n1982; //CHANX (4,2) #12 2002 2758 2741 1075
wire n1983; //CHANX (4,2) #13 1963 2660 2635 1075
wire n1984; //CHANX (4,2) #14 2004 2756 2743 1107
wire n1985; //CHANX (4,2) #15 1965 2662 2633 1107
wire n1986; //CHANX (4,2) #16 2006 2754 2745 1079
wire n1987; //CHANX (4,2) #17 1967 2664 2631 1079
wire n1988; //CHANX (4,2) #18 2008 2752 2747 1111
wire n1989; //CHANX (4,2) #19 1969 2666 2649 1111
wire n1990; //CHANX (5,2) #0 2850 2831 1349 1317
wire n1991; //CHANX (5,2) #1 1971 2768 2747 1349 1317
wire n1992; //CHANX (5,2) #2 2852 2833 1321
wire n1993; //CHANX (5,2) #3 1973 2750 2745 1321
wire n1994; //CHANX (5,2) #4 2854 2835 1353
wire n1995; //CHANX (5,2) #5 1975 2752 2743 1353
wire n1996; //CHANX (5,2) #6 2856 2837 1325
wire n1997; //CHANX (5,2) #7 1977 2754 2741 1325
wire n1998; //CHANX (5,2) #8 2858 2839 1357
wire n1999; //CHANX (5,2) #9 1979 2756 2739 1357
wire n2000; //CHANX (5,2) #10 2860 2841 1349 1317
wire n2001; //CHANX (5,2) #11 1981 2758 2737 1349 1317
wire n2002; //CHANX (5,2) #12 2862 2843 1321
wire n2003; //CHANX (5,2) #13 1983 2760 2735 1321
wire n2004; //CHANX (5,2) #14 2864 2845 1353
wire n2005; //CHANX (5,2) #15 1985 2762 2733 1353
wire n2006; //CHANX (5,2) #16 2866 2847 1325
wire n2007; //CHANX (5,2) #17 1987 2764 2731 1325
wire n2008; //CHANX (5,2) #18 2868 2849 1357
wire n2009; //CHANX (5,2) #19 1989 2766 2749 1357
wire n2010; //CHANX (1,3) #0 2030 2470 2469 395 363
wire n2011; //CHANX (1,3) #1 2370 2351 395 363
wire n2012; //CHANX (1,3) #2 2032 2488 2451 367
wire n2013; //CHANX (1,3) #3 2372 2353 367
wire n2014; //CHANX (1,3) #4 2034 2486 2453 399
wire n2015; //CHANX (1,3) #5 2374 2355 399
wire n2016; //CHANX (1,3) #6 2036 2484 2455 371
wire n2017; //CHANX (1,3) #7 2376 2357 371
wire n2018; //CHANX (1,3) #8 2038 2482 2457 403
wire n2019; //CHANX (1,3) #9 2378 2359 403
wire n2020; //CHANX (1,3) #10 2040 2480 2459 395 363
wire n2021; //CHANX (1,3) #11 2380 2361 395 363
wire n2022; //CHANX (1,3) #12 2042 2478 2461 367
wire n2023; //CHANX (1,3) #13 2382 2363 367
wire n2024; //CHANX (1,3) #14 2044 2476 2463 399
wire n2025; //CHANX (1,3) #15 2384 2365 399
wire n2026; //CHANX (1,3) #16 2046 2474 2465 371
wire n2027; //CHANX (1,3) #17 2386 2367 371
wire n2028; //CHANX (1,3) #18 2048 2472 2467 403
wire n2029; //CHANX (1,3) #19 2388 2369 403
wire n2030; //CHANX (2,3) #0 2050 2570 2569 641 609
wire n2031; //CHANX (2,3) #1 2011 2488 2467 641 609
wire n2032; //CHANX (2,3) #2 2052 2588 2551 613
wire n2033; //CHANX (2,3) #3 2013 2470 2465 613
wire n2034; //CHANX (2,3) #4 2054 2586 2553 645
wire n2035; //CHANX (2,3) #5 2015 2472 2463 645
wire n2036; //CHANX (2,3) #6 2056 2584 2555 617
wire n2037; //CHANX (2,3) #7 2017 2474 2461 617
wire n2038; //CHANX (2,3) #8 2058 2582 2557 649
wire n2039; //CHANX (2,3) #9 2019 2476 2459 649
wire n2040; //CHANX (2,3) #10 2060 2580 2559 641 609
wire n2041; //CHANX (2,3) #11 2021 2478 2457 641 609
wire n2042; //CHANX (2,3) #12 2062 2578 2561 613
wire n2043; //CHANX (2,3) #13 2023 2480 2455 613
wire n2044; //CHANX (2,3) #14 2064 2576 2563 645
wire n2045; //CHANX (2,3) #15 2025 2482 2453 645
wire n2046; //CHANX (2,3) #16 2066 2574 2565 617
wire n2047; //CHANX (2,3) #17 2027 2484 2451 617
wire n2048; //CHANX (2,3) #18 2068 2572 2567 649
wire n2049; //CHANX (2,3) #19 2029 2486 2469 649
wire n2050; //CHANX (3,3) #0 2070 2670 2669 887 855
wire n2051; //CHANX (3,3) #1 2031 2588 2567 887 855
wire n2052; //CHANX (3,3) #2 2072 2688 2651 859
wire n2053; //CHANX (3,3) #3 2033 2570 2565 859
wire n2054; //CHANX (3,3) #4 2074 2686 2653 891
wire n2055; //CHANX (3,3) #5 2035 2572 2563 891
wire n2056; //CHANX (3,3) #6 2076 2684 2655 863
wire n2057; //CHANX (3,3) #7 2037 2574 2561 863
wire n2058; //CHANX (3,3) #8 2078 2682 2657 895
wire n2059; //CHANX (3,3) #9 2039 2576 2559 895
wire n2060; //CHANX (3,3) #10 2080 2680 2659 887 855
wire n2061; //CHANX (3,3) #11 2041 2578 2557 887 855
wire n2062; //CHANX (3,3) #12 2082 2678 2661 859
wire n2063; //CHANX (3,3) #13 2043 2580 2555 859
wire n2064; //CHANX (3,3) #14 2084 2676 2663 891
wire n2065; //CHANX (3,3) #15 2045 2582 2553 891
wire n2066; //CHANX (3,3) #16 2086 2674 2665 863
wire n2067; //CHANX (3,3) #17 2047 2584 2551 863
wire n2068; //CHANX (3,3) #18 2088 2672 2667 895
wire n2069; //CHANX (3,3) #19 2049 2586 2569 895
wire n2070; //CHANX (4,3) #0 2090 2770 2769 1133 1101
wire n2071; //CHANX (4,3) #1 2051 2688 2667 1133 1101
wire n2072; //CHANX (4,3) #2 2092 2788 2751 1105
wire n2073; //CHANX (4,3) #3 2053 2670 2665 1105
wire n2074; //CHANX (4,3) #4 2094 2786 2753 1137
wire n2075; //CHANX (4,3) #5 2055 2672 2663 1137
wire n2076; //CHANX (4,3) #6 2096 2784 2755 1109
wire n2077; //CHANX (4,3) #7 2057 2674 2661 1109
wire n2078; //CHANX (4,3) #8 2098 2782 2757 1141
wire n2079; //CHANX (4,3) #9 2059 2676 2659 1141
wire n2080; //CHANX (4,3) #10 2100 2780 2759 1133 1101
wire n2081; //CHANX (4,3) #11 2061 2678 2657 1133 1101
wire n2082; //CHANX (4,3) #12 2102 2778 2761 1105
wire n2083; //CHANX (4,3) #13 2063 2680 2655 1105
wire n2084; //CHANX (4,3) #14 2104 2776 2763 1137
wire n2085; //CHANX (4,3) #15 2065 2682 2653 1137
wire n2086; //CHANX (4,3) #16 2106 2774 2765 1109
wire n2087; //CHANX (4,3) #17 2067 2684 2651 1109
wire n2088; //CHANX (4,3) #18 2108 2772 2767 1141
wire n2089; //CHANX (4,3) #19 2069 2686 2669 1141
wire n2090; //CHANX (5,3) #0 2870 2851 1379 1347
wire n2091; //CHANX (5,3) #1 2071 2788 2767 1379 1347
wire n2092; //CHANX (5,3) #2 2872 2853 1351
wire n2093; //CHANX (5,3) #3 2073 2770 2765 1351
wire n2094; //CHANX (5,3) #4 2874 2855 1383
wire n2095; //CHANX (5,3) #5 2075 2772 2763 1383
wire n2096; //CHANX (5,3) #6 2876 2857 1355
wire n2097; //CHANX (5,3) #7 2077 2774 2761 1355
wire n2098; //CHANX (5,3) #8 2878 2859 1387
wire n2099; //CHANX (5,3) #9 2079 2776 2759 1387
wire n2100; //CHANX (5,3) #10 2880 2861 1379 1347
wire n2101; //CHANX (5,3) #11 2081 2778 2757 1379 1347
wire n2102; //CHANX (5,3) #12 2882 2863 1351
wire n2103; //CHANX (5,3) #13 2083 2780 2755 1351
wire n2104; //CHANX (5,3) #14 2884 2865 1383
wire n2105; //CHANX (5,3) #15 2085 2782 2753 1383
wire n2106; //CHANX (5,3) #16 2886 2867 1355
wire n2107; //CHANX (5,3) #17 2087 2784 2751 1355
wire n2108; //CHANX (5,3) #18 2888 2869 1387
wire n2109; //CHANX (5,3) #19 2089 2786 2769 1387
wire n2110; //CHANX (1,4) #0 2130 2490 2489 425 393
wire n2111; //CHANX (1,4) #1 2390 2371 425 393
wire n2112; //CHANX (1,4) #2 2132 2508 2471 397
wire n2113; //CHANX (1,4) #3 2392 2373 397
wire n2114; //CHANX (1,4) #4 2134 2506 2473 429
wire n2115; //CHANX (1,4) #5 2394 2375 429
wire n2116; //CHANX (1,4) #6 2136 2504 2475 401
wire n2117; //CHANX (1,4) #7 2396 2377 401
wire n2118; //CHANX (1,4) #8 2138 2502 2477 433
wire n2119; //CHANX (1,4) #9 2398 2379 433
wire n2120; //CHANX (1,4) #10 2140 2500 2479 425 393
wire n2121; //CHANX (1,4) #11 2400 2381 425 393
wire n2122; //CHANX (1,4) #12 2142 2498 2481 397
wire n2123; //CHANX (1,4) #13 2402 2383 397
wire n2124; //CHANX (1,4) #14 2144 2496 2483 429
wire n2125; //CHANX (1,4) #15 2404 2385 429
wire n2126; //CHANX (1,4) #16 2146 2494 2485 401
wire n2127; //CHANX (1,4) #17 2406 2387 401
wire n2128; //CHANX (1,4) #18 2148 2492 2487 433
wire n2129; //CHANX (1,4) #19 2408 2389 433
wire n2130; //CHANX (2,4) #0 2150 2590 2589 671 639
wire n2131; //CHANX (2,4) #1 2111 2508 2487 671 639
wire n2132; //CHANX (2,4) #2 2152 2608 2571 643
wire n2133; //CHANX (2,4) #3 2113 2490 2485 643
wire n2134; //CHANX (2,4) #4 2154 2606 2573 675
wire n2135; //CHANX (2,4) #5 2115 2492 2483 675
wire n2136; //CHANX (2,4) #6 2156 2604 2575 647
wire n2137; //CHANX (2,4) #7 2117 2494 2481 647
wire n2138; //CHANX (2,4) #8 2158 2602 2577 679
wire n2139; //CHANX (2,4) #9 2119 2496 2479 679
wire n2140; //CHANX (2,4) #10 2160 2600 2579 671 639
wire n2141; //CHANX (2,4) #11 2121 2498 2477 671 639
wire n2142; //CHANX (2,4) #12 2162 2598 2581 643
wire n2143; //CHANX (2,4) #13 2123 2500 2475 643
wire n2144; //CHANX (2,4) #14 2164 2596 2583 675
wire n2145; //CHANX (2,4) #15 2125 2502 2473 675
wire n2146; //CHANX (2,4) #16 2166 2594 2585 647
wire n2147; //CHANX (2,4) #17 2127 2504 2471 647
wire n2148; //CHANX (2,4) #18 2168 2592 2587 679
wire n2149; //CHANX (2,4) #19 2129 2506 2489 679
wire n2150; //CHANX (3,4) #0 2170 2690 2689 917 885
wire n2151; //CHANX (3,4) #1 2131 2608 2587 917 885
wire n2152; //CHANX (3,4) #2 2172 2708 2671 889
wire n2153; //CHANX (3,4) #3 2133 2590 2585 889
wire n2154; //CHANX (3,4) #4 2174 2706 2673 921
wire n2155; //CHANX (3,4) #5 2135 2592 2583 921
wire n2156; //CHANX (3,4) #6 2176 2704 2675 893
wire n2157; //CHANX (3,4) #7 2137 2594 2581 893
wire n2158; //CHANX (3,4) #8 2178 2702 2677 925
wire n2159; //CHANX (3,4) #9 2139 2596 2579 925
wire n2160; //CHANX (3,4) #10 2180 2700 2679 917 885
wire n2161; //CHANX (3,4) #11 2141 2598 2577 917 885
wire n2162; //CHANX (3,4) #12 2182 2698 2681 889
wire n2163; //CHANX (3,4) #13 2143 2600 2575 889
wire n2164; //CHANX (3,4) #14 2184 2696 2683 921
wire n2165; //CHANX (3,4) #15 2145 2602 2573 921
wire n2166; //CHANX (3,4) #16 2186 2694 2685 893
wire n2167; //CHANX (3,4) #17 2147 2604 2571 893
wire n2168; //CHANX (3,4) #18 2188 2692 2687 925
wire n2169; //CHANX (3,4) #19 2149 2606 2589 925
wire n2170; //CHANX (4,4) #0 2190 2790 2789 1163 1131
wire n2171; //CHANX (4,4) #1 2151 2708 2687 1163 1131
wire n2172; //CHANX (4,4) #2 2192 2808 2771 1135
wire n2173; //CHANX (4,4) #3 2153 2690 2685 1135
wire n2174; //CHANX (4,4) #4 2194 2806 2773 1167
wire n2175; //CHANX (4,4) #5 2155 2692 2683 1167
wire n2176; //CHANX (4,4) #6 2196 2804 2775 1139
wire n2177; //CHANX (4,4) #7 2157 2694 2681 1139
wire n2178; //CHANX (4,4) #8 2198 2802 2777 1171
wire n2179; //CHANX (4,4) #9 2159 2696 2679 1171
wire n2180; //CHANX (4,4) #10 2200 2800 2779 1163 1131
wire n2181; //CHANX (4,4) #11 2161 2698 2677 1163 1131
wire n2182; //CHANX (4,4) #12 2202 2798 2781 1135
wire n2183; //CHANX (4,4) #13 2163 2700 2675 1135
wire n2184; //CHANX (4,4) #14 2204 2796 2783 1167
wire n2185; //CHANX (4,4) #15 2165 2702 2673 1167
wire n2186; //CHANX (4,4) #16 2206 2794 2785 1139
wire n2187; //CHANX (4,4) #17 2167 2704 2671 1139
wire n2188; //CHANX (4,4) #18 2208 2792 2787 1171
wire n2189; //CHANX (4,4) #19 2169 2706 2689 1171
wire n2190; //CHANX (5,4) #0 2890 2871 1409 1377
wire n2191; //CHANX (5,4) #1 2171 2808 2787 1409 1377
wire n2192; //CHANX (5,4) #2 2892 2873 1381
wire n2193; //CHANX (5,4) #3 2173 2790 2785 1381
wire n2194; //CHANX (5,4) #4 2894 2875 1413
wire n2195; //CHANX (5,4) #5 2175 2792 2783 1413
wire n2196; //CHANX (5,4) #6 2896 2877 1385
wire n2197; //CHANX (5,4) #7 2177 2794 2781 1385
wire n2198; //CHANX (5,4) #8 2898 2879 1417
wire n2199; //CHANX (5,4) #9 2179 2796 2779 1417
wire n2200; //CHANX (5,4) #10 2900 2881 1409 1377
wire n2201; //CHANX (5,4) #11 2181 2798 2777 1409 1377
wire n2202; //CHANX (5,4) #12 2902 2883 1381
wire n2203; //CHANX (5,4) #13 2183 2800 2775 1381
wire n2204; //CHANX (5,4) #14 2904 2885 1413
wire n2205; //CHANX (5,4) #15 2185 2802 2773 1413
wire n2206; //CHANX (5,4) #16 2906 2887 1385
wire n2207; //CHANX (5,4) #17 2187 2804 2771 1385
wire n2208; //CHANX (5,4) #18 2908 2889 1417
wire n2209; //CHANX (5,4) #19 2189 2806 2789 1417
wire n2210; //CHANX (1,5) #0 2230 2491 465 462 423
wire n2211; //CHANX (1,5) #1 2407 465 462 423
wire n2212; //CHANX (1,5) #2 2232 2497 468 427
wire n2213; //CHANX (1,5) #3 2405 468 427
wire n2214; //CHANX (1,5) #4 2234 2503 474 471
wire n2215; //CHANX (1,5) #5 2403 474 471
wire n2216; //CHANX (1,5) #6 2236 2509 477 431
wire n2217; //CHANX (1,5) #7 2401 477 431
wire n2218; //CHANX (1,5) #8 2238 2493 483 480
wire n2219; //CHANX (1,5) #9 2399 483 480
wire n2220; //CHANX (1,5) #10 2240 2495 465 462 423
wire n2221; //CHANX (1,5) #11 2397 465 462 423
wire n2222; //CHANX (1,5) #12 2242 2499 468 427
wire n2223; //CHANX (1,5) #13 2395 468 427
wire n2224; //CHANX (1,5) #14 2244 2501 474 471
wire n2225; //CHANX (1,5) #15 2393 474 471
wire n2226; //CHANX (1,5) #16 2246 2505 477 431
wire n2227; //CHANX (1,5) #17 2391 477 431
wire n2228; //CHANX (1,5) #18 2248 2507 483 480
wire n2229; //CHANX (1,5) #19 2409 483 480
wire n2230; //CHANX (2,5) #0 2250 2591 711 708 669
wire n2231; //CHANX (2,5) #1 2211 2491 711 708 669
wire n2232; //CHANX (2,5) #2 2252 2597 714 673
wire n2233; //CHANX (2,5) #3 2213 2497 714 673
wire n2234; //CHANX (2,5) #4 2254 2603 720 717
wire n2235; //CHANX (2,5) #5 2215 2503 720 717
wire n2236; //CHANX (2,5) #6 2256 2609 723 677
wire n2237; //CHANX (2,5) #7 2217 2509 723 677
wire n2238; //CHANX (2,5) #8 2258 2593 729 726
wire n2239; //CHANX (2,5) #9 2219 2493 729 726
wire n2240; //CHANX (2,5) #10 2260 2595 711 708 669
wire n2241; //CHANX (2,5) #11 2221 2495 711 708 669
wire n2242; //CHANX (2,5) #12 2262 2599 714 673
wire n2243; //CHANX (2,5) #13 2223 2499 714 673
wire n2244; //CHANX (2,5) #14 2264 2601 720 717
wire n2245; //CHANX (2,5) #15 2225 2501 720 717
wire n2246; //CHANX (2,5) #16 2266 2605 723 677
wire n2247; //CHANX (2,5) #17 2227 2505 723 677
wire n2248; //CHANX (2,5) #18 2268 2607 729 726
wire n2249; //CHANX (2,5) #19 2229 2507 729 726
wire n2250; //CHANX (3,5) #0 2270 2691 957 954 915
wire n2251; //CHANX (3,5) #1 2231 2591 957 954 915
wire n2252; //CHANX (3,5) #2 2272 2697 960 919
wire n2253; //CHANX (3,5) #3 2233 2597 960 919
wire n2254; //CHANX (3,5) #4 2274 2703 966 963
wire n2255; //CHANX (3,5) #5 2235 2603 966 963
wire n2256; //CHANX (3,5) #6 2276 2709 969 923
wire n2257; //CHANX (3,5) #7 2237 2609 969 923
wire n2258; //CHANX (3,5) #8 2278 2693 975 972
wire n2259; //CHANX (3,5) #9 2239 2593 975 972
wire n2260; //CHANX (3,5) #10 2280 2695 957 954 915
wire n2261; //CHANX (3,5) #11 2241 2595 957 954 915
wire n2262; //CHANX (3,5) #12 2282 2699 960 919
wire n2263; //CHANX (3,5) #13 2243 2599 960 919
wire n2264; //CHANX (3,5) #14 2284 2701 966 963
wire n2265; //CHANX (3,5) #15 2245 2601 966 963
wire n2266; //CHANX (3,5) #16 2286 2705 969 923
wire n2267; //CHANX (3,5) #17 2247 2605 969 923
wire n2268; //CHANX (3,5) #18 2288 2707 975 972
wire n2269; //CHANX (3,5) #19 2249 2607 975 972
wire n2270; //CHANX (4,5) #0 2290 2791 1203 1200 1161
wire n2271; //CHANX (4,5) #1 2251 2691 1203 1200 1161
wire n2272; //CHANX (4,5) #2 2292 2797 1206 1165
wire n2273; //CHANX (4,5) #3 2253 2697 1206 1165
wire n2274; //CHANX (4,5) #4 2294 2803 1212 1209
wire n2275; //CHANX (4,5) #5 2255 2703 1212 1209
wire n2276; //CHANX (4,5) #6 2296 2809 1215 1169
wire n2277; //CHANX (4,5) #7 2257 2709 1215 1169
wire n2278; //CHANX (4,5) #8 2298 2793 1221 1218
wire n2279; //CHANX (4,5) #9 2259 2693 1221 1218
wire n2280; //CHANX (4,5) #10 2300 2795 1203 1200 1161
wire n2281; //CHANX (4,5) #11 2261 2695 1203 1200 1161
wire n2282; //CHANX (4,5) #12 2302 2799 1206 1165
wire n2283; //CHANX (4,5) #13 2263 2699 1206 1165
wire n2284; //CHANX (4,5) #14 2304 2801 1212 1209
wire n2285; //CHANX (4,5) #15 2265 2701 1212 1209
wire n2286; //CHANX (4,5) #16 2306 2805 1215 1169
wire n2287; //CHANX (4,5) #17 2267 2705 1215 1169
wire n2288; //CHANX (4,5) #18 2308 2807 1221 1218
wire n2289; //CHANX (4,5) #19 2269 2707 1221 1218
wire n2290; //CHANX (5,5) #0 2909 1449 1446 1407
wire n2291; //CHANX (5,5) #1 2271 2791 1449 1446 1407
wire n2292; //CHANX (5,5) #2 2891 1452 1411
wire n2293; //CHANX (5,5) #3 2273 2797 1452 1411
wire n2294; //CHANX (5,5) #4 2893 1458 1455
wire n2295; //CHANX (5,5) #5 2275 2803 1458 1455
wire n2296; //CHANX (5,5) #6 2895 1461 1415
wire n2297; //CHANX (5,5) #7 2277 2809 1461 1415
wire n2298; //CHANX (5,5) #8 2897 1467 1464
wire n2299; //CHANX (5,5) #9 2279 2793 1467 1464
wire n2300; //CHANX (5,5) #10 2899 1449 1446 1407
wire n2301; //CHANX (5,5) #11 2281 2795 1449 1446 1407
wire n2302; //CHANX (5,5) #12 2901 1452 1411
wire n2303; //CHANX (5,5) #13 2283 2799 1452 1411
wire n2304; //CHANX (5,5) #14 2903 1458 1455
wire n2305; //CHANX (5,5) #15 2285 2801 1458 1455
wire n2306; //CHANX (5,5) #16 2905 1461 1415
wire n2307; //CHANX (5,5) #17 2287 2805 1461 1415
wire n2308; //CHANX (5,5) #18 2907 1467 1464
wire n2309; //CHANX (5,5) #19 2289 2807 1467 1464
wire n2310; //CHANY (0,1) #0 2330 1814 27 24
wire n2311; //CHANY (0,1) #1 1712 27 24
wire n2312; //CHANY (0,1) #2 2332 1820 306 30
wire n2313; //CHANY (0,1) #3 1714 306 30
wire n2314; //CHANY (0,1) #4 2334 1826 310 36 33
wire n2315; //CHANY (0,1) #5 1716 310 36 33
wire n2316; //CHANY (0,1) #6 2336 1810 42 39
wire n2317; //CHANY (0,1) #7 1718 42 39
wire n2318; //CHANY (0,1) #8 2338 1812 314 45
wire n2319; //CHANY (0,1) #9 1720 314 45
wire n2320; //CHANY (0,1) #10 2340 1816 27 24
wire n2321; //CHANY (0,1) #11 1722 27 24
wire n2322; //CHANY (0,1) #12 2342 1818 306 30
wire n2323; //CHANY (0,1) #13 1724 306 30
wire n2324; //CHANY (0,1) #14 2344 1822 310 36 33
wire n2325; //CHANY (0,1) #15 1726 310 36 33
wire n2326; //CHANY (0,1) #16 2346 1824 42 39
wire n2327; //CHANY (0,1) #17 1728 42 39
wire n2328; //CHANY (0,1) #18 2348 1828 314 45
wire n2329; //CHANY (0,1) #19 1710 314 45
wire n2330; //CHANY (0,2) #0 2350 1914 75 72
wire n2331; //CHANY (0,2) #1 2311 1814 75 72
wire n2332; //CHANY (0,2) #2 2352 1920 336 78
wire n2333; //CHANY (0,2) #3 2313 1820 336 78
wire n2334; //CHANY (0,2) #4 2354 1926 340 84 81
wire n2335; //CHANY (0,2) #5 2315 1826 340 84 81
wire n2336; //CHANY (0,2) #6 2356 1910 90 87
wire n2337; //CHANY (0,2) #7 2317 1810 90 87
wire n2338; //CHANY (0,2) #8 2358 1912 344 93
wire n2339; //CHANY (0,2) #9 2319 1812 344 93
wire n2340; //CHANY (0,2) #10 2360 1916 75 72
wire n2341; //CHANY (0,2) #11 2321 1816 75 72
wire n2342; //CHANY (0,2) #12 2362 1918 336 78
wire n2343; //CHANY (0,2) #13 2323 1818 336 78
wire n2344; //CHANY (0,2) #14 2364 1922 340 84 81
wire n2345; //CHANY (0,2) #15 2325 1822 340 84 81
wire n2346; //CHANY (0,2) #16 2366 1924 90 87
wire n2347; //CHANY (0,2) #17 2327 1824 90 87
wire n2348; //CHANY (0,2) #18 2368 1928 344 93
wire n2349; //CHANY (0,2) #19 2329 1828 344 93
wire n2350; //CHANY (0,3) #0 2370 2014 123 120
wire n2351; //CHANY (0,3) #1 2331 1914 123 120
wire n2352; //CHANY (0,3) #2 2372 2020 366 126
wire n2353; //CHANY (0,3) #3 2333 1920 366 126
wire n2354; //CHANY (0,3) #4 2374 2026 370 132 129
wire n2355; //CHANY (0,3) #5 2335 1926 370 132 129
wire n2356; //CHANY (0,3) #6 2376 2010 138 135
wire n2357; //CHANY (0,3) #7 2337 1910 138 135
wire n2358; //CHANY (0,3) #8 2378 2012 374 141
wire n2359; //CHANY (0,3) #9 2339 1912 374 141
wire n2360; //CHANY (0,3) #10 2380 2016 123 120
wire n2361; //CHANY (0,3) #11 2341 1916 123 120
wire n2362; //CHANY (0,3) #12 2382 2018 366 126
wire n2363; //CHANY (0,3) #13 2343 1918 366 126
wire n2364; //CHANY (0,3) #14 2384 2022 370 132 129
wire n2365; //CHANY (0,3) #15 2345 1922 370 132 129
wire n2366; //CHANY (0,3) #16 2386 2024 138 135
wire n2367; //CHANY (0,3) #17 2347 1924 138 135
wire n2368; //CHANY (0,3) #18 2388 2028 374 141
wire n2369; //CHANY (0,3) #19 2349 1928 374 141
wire n2370; //CHANY (0,4) #0 2390 2114 171 168
wire n2371; //CHANY (0,4) #1 2351 2014 171 168
wire n2372; //CHANY (0,4) #2 2392 2120 396 174
wire n2373; //CHANY (0,4) #3 2353 2020 396 174
wire n2374; //CHANY (0,4) #4 2394 2126 400 180 177
wire n2375; //CHANY (0,4) #5 2355 2026 400 180 177
wire n2376; //CHANY (0,4) #6 2396 2110 186 183
wire n2377; //CHANY (0,4) #7 2357 2010 186 183
wire n2378; //CHANY (0,4) #8 2398 2112 404 189
wire n2379; //CHANY (0,4) #9 2359 2012 404 189
wire n2380; //CHANY (0,4) #10 2400 2116 171 168
wire n2381; //CHANY (0,4) #11 2361 2016 171 168
wire n2382; //CHANY (0,4) #12 2402 2118 396 174
wire n2383; //CHANY (0,4) #13 2363 2018 396 174
wire n2384; //CHANY (0,4) #14 2404 2122 400 180 177
wire n2385; //CHANY (0,4) #15 2365 2022 400 180 177
wire n2386; //CHANY (0,4) #16 2406 2124 186 183
wire n2387; //CHANY (0,4) #17 2367 2024 186 183
wire n2388; //CHANY (0,4) #18 2408 2128 404 189
wire n2389; //CHANY (0,4) #19 2369 2028 404 189
wire n2390; //CHANY (0,5) #0 2226 219 216
wire n2391; //CHANY (0,5) #1 2371 2114 219 216
wire n2392; //CHANY (0,5) #2 2224 426 222
wire n2393; //CHANY (0,5) #3 2373 2120 426 222
wire n2394; //CHANY (0,5) #4 2222 430 228 225
wire n2395; //CHANY (0,5) #5 2375 2126 430 228 225
wire n2396; //CHANY (0,5) #6 2220 234 231
wire n2397; //CHANY (0,5) #7 2377 2110 234 231
wire n2398; //CHANY (0,5) #8 2218 434 237
wire n2399; //CHANY (0,5) #9 2379 2112 434 237
wire n2400; //CHANY (0,5) #10 2216 219 216
wire n2401; //CHANY (0,5) #11 2381 2116 219 216
wire n2402; //CHANY (0,5) #12 2214 426 222
wire n2403; //CHANY (0,5) #13 2383 2118 426 222
wire n2404; //CHANY (0,5) #14 2212 430 228 225
wire n2405; //CHANY (0,5) #15 2385 2122 430 228 225
wire n2406; //CHANY (0,5) #16 2210 234 231
wire n2407; //CHANY (0,5) #17 2387 2124 234 231
wire n2408; //CHANY (0,5) #18 2228 434 237
wire n2409; //CHANY (0,5) #19 2389 2128 434 237
wire n2410; //CHANY (1,1) #0 2430 1846 1813 304
wire n2411; //CHANY (1,1) #1 1730 1711 304
wire n2412; //CHANY (1,1) #2 2432 1844 1815 552
wire n2413; //CHANY (1,1) #3 1732 1713 552
wire n2414; //CHANY (1,1) #4 2434 1842 1817 556 308
wire n2415; //CHANY (1,1) #5 1734 1715 556 308
wire n2416; //CHANY (1,1) #6 2436 1840 1819 312
wire n2417; //CHANY (1,1) #7 1736 1717 312
wire n2418; //CHANY (1,1) #8 2438 1838 1821 560
wire n2419; //CHANY (1,1) #9 1738 1719 560
wire n2420; //CHANY (1,1) #10 2440 1836 1823 304
wire n2421; //CHANY (1,1) #11 1740 1721 304
wire n2422; //CHANY (1,1) #12 2442 1834 1825 552
wire n2423; //CHANY (1,1) #13 1742 1723 552
wire n2424; //CHANY (1,1) #14 2444 1832 1827 556 308
wire n2425; //CHANY (1,1) #15 1744 1725 556 308
wire n2426; //CHANY (1,1) #16 2446 1830 1829 312
wire n2427; //CHANY (1,1) #17 1746 1727 312
wire n2428; //CHANY (1,1) #18 2448 1848 1811 560
wire n2429; //CHANY (1,1) #19 1748 1729 560
wire n2430; //CHANY (1,2) #0 2450 1946 1913 334
wire n2431; //CHANY (1,2) #1 2411 1832 1811 334
wire n2432; //CHANY (1,2) #2 2452 1944 1915 582
wire n2433; //CHANY (1,2) #3 2413 1834 1829 582
wire n2434; //CHANY (1,2) #4 2454 1942 1917 586 338
wire n2435; //CHANY (1,2) #5 2415 1836 1827 586 338
wire n2436; //CHANY (1,2) #6 2456 1940 1919 342
wire n2437; //CHANY (1,2) #7 2417 1838 1825 342
wire n2438; //CHANY (1,2) #8 2458 1938 1921 590
wire n2439; //CHANY (1,2) #9 2419 1840 1823 590
wire n2440; //CHANY (1,2) #10 2460 1936 1923 334
wire n2441; //CHANY (1,2) #11 2421 1842 1821 334
wire n2442; //CHANY (1,2) #12 2462 1934 1925 582
wire n2443; //CHANY (1,2) #13 2423 1844 1819 582
wire n2444; //CHANY (1,2) #14 2464 1932 1927 586 338
wire n2445; //CHANY (1,2) #15 2425 1846 1817 586 338
wire n2446; //CHANY (1,2) #16 2466 1930 1929 342
wire n2447; //CHANY (1,2) #17 2427 1848 1815 342
wire n2448; //CHANY (1,2) #18 2468 1948 1911 590
wire n2449; //CHANY (1,2) #19 2429 1830 1813 590
wire n2450; //CHANY (1,3) #0 2470 2046 2013 364
wire n2451; //CHANY (1,3) #1 2431 1932 1911 364
wire n2452; //CHANY (1,3) #2 2472 2044 2015 612
wire n2453; //CHANY (1,3) #3 2433 1934 1929 612
wire n2454; //CHANY (1,3) #4 2474 2042 2017 616 368
wire n2455; //CHANY (1,3) #5 2435 1936 1927 616 368
wire n2456; //CHANY (1,3) #6 2476 2040 2019 372
wire n2457; //CHANY (1,3) #7 2437 1938 1925 372
wire n2458; //CHANY (1,3) #8 2478 2038 2021 620
wire n2459; //CHANY (1,3) #9 2439 1940 1923 620
wire n2460; //CHANY (1,3) #10 2480 2036 2023 364
wire n2461; //CHANY (1,3) #11 2441 1942 1921 364
wire n2462; //CHANY (1,3) #12 2482 2034 2025 612
wire n2463; //CHANY (1,3) #13 2443 1944 1919 612
wire n2464; //CHANY (1,3) #14 2484 2032 2027 616 368
wire n2465; //CHANY (1,3) #15 2445 1946 1917 616 368
wire n2466; //CHANY (1,3) #16 2486 2030 2029 372
wire n2467; //CHANY (1,3) #17 2447 1948 1915 372
wire n2468; //CHANY (1,3) #18 2488 2048 2011 620
wire n2469; //CHANY (1,3) #19 2449 1930 1913 620
wire n2470; //CHANY (1,4) #0 2490 2146 2113 394
wire n2471; //CHANY (1,4) #1 2451 2032 2011 394
wire n2472; //CHANY (1,4) #2 2492 2144 2115 642
wire n2473; //CHANY (1,4) #3 2453 2034 2029 642
wire n2474; //CHANY (1,4) #4 2494 2142 2117 646 398
wire n2475; //CHANY (1,4) #5 2455 2036 2027 646 398
wire n2476; //CHANY (1,4) #6 2496 2140 2119 402
wire n2477; //CHANY (1,4) #7 2457 2038 2025 402
wire n2478; //CHANY (1,4) #8 2498 2138 2121 650
wire n2479; //CHANY (1,4) #9 2459 2040 2023 650
wire n2480; //CHANY (1,4) #10 2500 2136 2123 394
wire n2481; //CHANY (1,4) #11 2461 2042 2021 394
wire n2482; //CHANY (1,4) #12 2502 2134 2125 642
wire n2483; //CHANY (1,4) #13 2463 2044 2019 642
wire n2484; //CHANY (1,4) #14 2504 2132 2127 646 398
wire n2485; //CHANY (1,4) #15 2465 2046 2017 646 398
wire n2486; //CHANY (1,4) #16 2506 2130 2129 402
wire n2487; //CHANY (1,4) #17 2467 2048 2015 402
wire n2488; //CHANY (1,4) #18 2508 2148 2111 650
wire n2489; //CHANY (1,4) #19 2469 2030 2013 650
wire n2490; //CHANY (1,5) #0 2230 2211 424
wire n2491; //CHANY (1,5) #1 2471 2132 2111 424
wire n2492; //CHANY (1,5) #2 2232 2213 672
wire n2493; //CHANY (1,5) #3 2473 2134 2129 672
wire n2494; //CHANY (1,5) #4 2234 2215 676 428
wire n2495; //CHANY (1,5) #5 2475 2136 2127 676 428
wire n2496; //CHANY (1,5) #6 2236 2217 432
wire n2497; //CHANY (1,5) #7 2477 2138 2125 432
wire n2498; //CHANY (1,5) #8 2238 2219 680
wire n2499; //CHANY (1,5) #9 2479 2140 2123 680
wire n2500; //CHANY (1,5) #10 2240 2221 424
wire n2501; //CHANY (1,5) #11 2481 2142 2121 424
wire n2502; //CHANY (1,5) #12 2242 2223 672
wire n2503; //CHANY (1,5) #13 2483 2144 2119 672
wire n2504; //CHANY (1,5) #14 2244 2225 676 428
wire n2505; //CHANY (1,5) #15 2485 2146 2117 676 428
wire n2506; //CHANY (1,5) #16 2246 2227 432
wire n2507; //CHANY (1,5) #17 2487 2148 2115 432
wire n2508; //CHANY (1,5) #18 2248 2229 680
wire n2509; //CHANY (1,5) #19 2489 2130 2113 680
wire n2510; //CHANY (2,1) #0 2530 1866 1833 550
wire n2511; //CHANY (2,1) #1 1750 1731 550
wire n2512; //CHANY (2,1) #2 2532 1864 1835 798
wire n2513; //CHANY (2,1) #3 1752 1733 798
wire n2514; //CHANY (2,1) #4 2534 1862 1837 802 554
wire n2515; //CHANY (2,1) #5 1754 1735 802 554
wire n2516; //CHANY (2,1) #6 2536 1860 1839 558
wire n2517; //CHANY (2,1) #7 1756 1737 558
wire n2518; //CHANY (2,1) #8 2538 1858 1841 806
wire n2519; //CHANY (2,1) #9 1758 1739 806
wire n2520; //CHANY (2,1) #10 2540 1856 1843 550
wire n2521; //CHANY (2,1) #11 1760 1741 550
wire n2522; //CHANY (2,1) #12 2542 1854 1845 798
wire n2523; //CHANY (2,1) #13 1762 1743 798
wire n2524; //CHANY (2,1) #14 2544 1852 1847 802 554
wire n2525; //CHANY (2,1) #15 1764 1745 802 554
wire n2526; //CHANY (2,1) #16 2546 1850 1849 558
wire n2527; //CHANY (2,1) #17 1766 1747 558
wire n2528; //CHANY (2,1) #18 2548 1868 1831 806
wire n2529; //CHANY (2,1) #19 1768 1749 806
wire n2530; //CHANY (2,2) #0 2550 1966 1933 580
wire n2531; //CHANY (2,2) #1 2511 1852 1831 580
wire n2532; //CHANY (2,2) #2 2552 1964 1935 828
wire n2533; //CHANY (2,2) #3 2513 1854 1849 828
wire n2534; //CHANY (2,2) #4 2554 1962 1937 832 584
wire n2535; //CHANY (2,2) #5 2515 1856 1847 832 584
wire n2536; //CHANY (2,2) #6 2556 1960 1939 588
wire n2537; //CHANY (2,2) #7 2517 1858 1845 588
wire n2538; //CHANY (2,2) #8 2558 1958 1941 836
wire n2539; //CHANY (2,2) #9 2519 1860 1843 836
wire n2540; //CHANY (2,2) #10 2560 1956 1943 580
wire n2541; //CHANY (2,2) #11 2521 1862 1841 580
wire n2542; //CHANY (2,2) #12 2562 1954 1945 828
wire n2543; //CHANY (2,2) #13 2523 1864 1839 828
wire n2544; //CHANY (2,2) #14 2564 1952 1947 832 584
wire n2545; //CHANY (2,2) #15 2525 1866 1837 832 584
wire n2546; //CHANY (2,2) #16 2566 1950 1949 588
wire n2547; //CHANY (2,2) #17 2527 1868 1835 588
wire n2548; //CHANY (2,2) #18 2568 1968 1931 836
wire n2549; //CHANY (2,2) #19 2529 1850 1833 836
wire n2550; //CHANY (2,3) #0 2570 2066 2033 610
wire n2551; //CHANY (2,3) #1 2531 1952 1931 610
wire n2552; //CHANY (2,3) #2 2572 2064 2035 858
wire n2553; //CHANY (2,3) #3 2533 1954 1949 858
wire n2554; //CHANY (2,3) #4 2574 2062 2037 862 614
wire n2555; //CHANY (2,3) #5 2535 1956 1947 862 614
wire n2556; //CHANY (2,3) #6 2576 2060 2039 618
wire n2557; //CHANY (2,3) #7 2537 1958 1945 618
wire n2558; //CHANY (2,3) #8 2578 2058 2041 866
wire n2559; //CHANY (2,3) #9 2539 1960 1943 866
wire n2560; //CHANY (2,3) #10 2580 2056 2043 610
wire n2561; //CHANY (2,3) #11 2541 1962 1941 610
wire n2562; //CHANY (2,3) #12 2582 2054 2045 858
wire n2563; //CHANY (2,3) #13 2543 1964 1939 858
wire n2564; //CHANY (2,3) #14 2584 2052 2047 862 614
wire n2565; //CHANY (2,3) #15 2545 1966 1937 862 614
wire n2566; //CHANY (2,3) #16 2586 2050 2049 618
wire n2567; //CHANY (2,3) #17 2547 1968 1935 618
wire n2568; //CHANY (2,3) #18 2588 2068 2031 866
wire n2569; //CHANY (2,3) #19 2549 1950 1933 866
wire n2570; //CHANY (2,4) #0 2590 2166 2133 640
wire n2571; //CHANY (2,4) #1 2551 2052 2031 640
wire n2572; //CHANY (2,4) #2 2592 2164 2135 888
wire n2573; //CHANY (2,4) #3 2553 2054 2049 888
wire n2574; //CHANY (2,4) #4 2594 2162 2137 892 644
wire n2575; //CHANY (2,4) #5 2555 2056 2047 892 644
wire n2576; //CHANY (2,4) #6 2596 2160 2139 648
wire n2577; //CHANY (2,4) #7 2557 2058 2045 648
wire n2578; //CHANY (2,4) #8 2598 2158 2141 896
wire n2579; //CHANY (2,4) #9 2559 2060 2043 896
wire n2580; //CHANY (2,4) #10 2600 2156 2143 640
wire n2581; //CHANY (2,4) #11 2561 2062 2041 640
wire n2582; //CHANY (2,4) #12 2602 2154 2145 888
wire n2583; //CHANY (2,4) #13 2563 2064 2039 888
wire n2584; //CHANY (2,4) #14 2604 2152 2147 892 644
wire n2585; //CHANY (2,4) #15 2565 2066 2037 892 644
wire n2586; //CHANY (2,4) #16 2606 2150 2149 648
wire n2587; //CHANY (2,4) #17 2567 2068 2035 648
wire n2588; //CHANY (2,4) #18 2608 2168 2131 896
wire n2589; //CHANY (2,4) #19 2569 2050 2033 896
wire n2590; //CHANY (2,5) #0 2250 2231 670
wire n2591; //CHANY (2,5) #1 2571 2152 2131 670
wire n2592; //CHANY (2,5) #2 2252 2233 918
wire n2593; //CHANY (2,5) #3 2573 2154 2149 918
wire n2594; //CHANY (2,5) #4 2254 2235 922 674
wire n2595; //CHANY (2,5) #5 2575 2156 2147 922 674
wire n2596; //CHANY (2,5) #6 2256 2237 678
wire n2597; //CHANY (2,5) #7 2577 2158 2145 678
wire n2598; //CHANY (2,5) #8 2258 2239 926
wire n2599; //CHANY (2,5) #9 2579 2160 2143 926
wire n2600; //CHANY (2,5) #10 2260 2241 670
wire n2601; //CHANY (2,5) #11 2581 2162 2141 670
wire n2602; //CHANY (2,5) #12 2262 2243 918
wire n2603; //CHANY (2,5) #13 2583 2164 2139 918
wire n2604; //CHANY (2,5) #14 2264 2245 922 674
wire n2605; //CHANY (2,5) #15 2585 2166 2137 922 674
wire n2606; //CHANY (2,5) #16 2266 2247 678
wire n2607; //CHANY (2,5) #17 2587 2168 2135 678
wire n2608; //CHANY (2,5) #18 2268 2249 926
wire n2609; //CHANY (2,5) #19 2589 2150 2133 926
wire n2610; //CHANY (3,1) #0 2630 1886 1853 796
wire n2611; //CHANY (3,1) #1 1770 1751 796
wire n2612; //CHANY (3,1) #2 2632 1884 1855 1044
wire n2613; //CHANY (3,1) #3 1772 1753 1044
wire n2614; //CHANY (3,1) #4 2634 1882 1857 1048 800
wire n2615; //CHANY (3,1) #5 1774 1755 1048 800
wire n2616; //CHANY (3,1) #6 2636 1880 1859 804
wire n2617; //CHANY (3,1) #7 1776 1757 804
wire n2618; //CHANY (3,1) #8 2638 1878 1861 1052
wire n2619; //CHANY (3,1) #9 1778 1759 1052
wire n2620; //CHANY (3,1) #10 2640 1876 1863 796
wire n2621; //CHANY (3,1) #11 1780 1761 796
wire n2622; //CHANY (3,1) #12 2642 1874 1865 1044
wire n2623; //CHANY (3,1) #13 1782 1763 1044
wire n2624; //CHANY (3,1) #14 2644 1872 1867 1048 800
wire n2625; //CHANY (3,1) #15 1784 1765 1048 800
wire n2626; //CHANY (3,1) #16 2646 1870 1869 804
wire n2627; //CHANY (3,1) #17 1786 1767 804
wire n2628; //CHANY (3,1) #18 2648 1888 1851 1052
wire n2629; //CHANY (3,1) #19 1788 1769 1052
wire n2630; //CHANY (3,2) #0 2650 1986 1953 826
wire n2631; //CHANY (3,2) #1 2611 1872 1851 826
wire n2632; //CHANY (3,2) #2 2652 1984 1955 1074
wire n2633; //CHANY (3,2) #3 2613 1874 1869 1074
wire n2634; //CHANY (3,2) #4 2654 1982 1957 1078 830
wire n2635; //CHANY (3,2) #5 2615 1876 1867 1078 830
wire n2636; //CHANY (3,2) #6 2656 1980 1959 834
wire n2637; //CHANY (3,2) #7 2617 1878 1865 834
wire n2638; //CHANY (3,2) #8 2658 1978 1961 1082
wire n2639; //CHANY (3,2) #9 2619 1880 1863 1082
wire n2640; //CHANY (3,2) #10 2660 1976 1963 826
wire n2641; //CHANY (3,2) #11 2621 1882 1861 826
wire n2642; //CHANY (3,2) #12 2662 1974 1965 1074
wire n2643; //CHANY (3,2) #13 2623 1884 1859 1074
wire n2644; //CHANY (3,2) #14 2664 1972 1967 1078 830
wire n2645; //CHANY (3,2) #15 2625 1886 1857 1078 830
wire n2646; //CHANY (3,2) #16 2666 1970 1969 834
wire n2647; //CHANY (3,2) #17 2627 1888 1855 834
wire n2648; //CHANY (3,2) #18 2668 1988 1951 1082
wire n2649; //CHANY (3,2) #19 2629 1870 1853 1082
wire n2650; //CHANY (3,3) #0 2670 2086 2053 856
wire n2651; //CHANY (3,3) #1 2631 1972 1951 856
wire n2652; //CHANY (3,3) #2 2672 2084 2055 1104
wire n2653; //CHANY (3,3) #3 2633 1974 1969 1104
wire n2654; //CHANY (3,3) #4 2674 2082 2057 1108 860
wire n2655; //CHANY (3,3) #5 2635 1976 1967 1108 860
wire n2656; //CHANY (3,3) #6 2676 2080 2059 864
wire n2657; //CHANY (3,3) #7 2637 1978 1965 864
wire n2658; //CHANY (3,3) #8 2678 2078 2061 1112
wire n2659; //CHANY (3,3) #9 2639 1980 1963 1112
wire n2660; //CHANY (3,3) #10 2680 2076 2063 856
wire n2661; //CHANY (3,3) #11 2641 1982 1961 856
wire n2662; //CHANY (3,3) #12 2682 2074 2065 1104
wire n2663; //CHANY (3,3) #13 2643 1984 1959 1104
wire n2664; //CHANY (3,3) #14 2684 2072 2067 1108 860
wire n2665; //CHANY (3,3) #15 2645 1986 1957 1108 860
wire n2666; //CHANY (3,3) #16 2686 2070 2069 864
wire n2667; //CHANY (3,3) #17 2647 1988 1955 864
wire n2668; //CHANY (3,3) #18 2688 2088 2051 1112
wire n2669; //CHANY (3,3) #19 2649 1970 1953 1112
wire n2670; //CHANY (3,4) #0 2690 2186 2153 886
wire n2671; //CHANY (3,4) #1 2651 2072 2051 886
wire n2672; //CHANY (3,4) #2 2692 2184 2155 1134
wire n2673; //CHANY (3,4) #3 2653 2074 2069 1134
wire n2674; //CHANY (3,4) #4 2694 2182 2157 1138 890
wire n2675; //CHANY (3,4) #5 2655 2076 2067 1138 890
wire n2676; //CHANY (3,4) #6 2696 2180 2159 894
wire n2677; //CHANY (3,4) #7 2657 2078 2065 894
wire n2678; //CHANY (3,4) #8 2698 2178 2161 1142
wire n2679; //CHANY (3,4) #9 2659 2080 2063 1142
wire n2680; //CHANY (3,4) #10 2700 2176 2163 886
wire n2681; //CHANY (3,4) #11 2661 2082 2061 886
wire n2682; //CHANY (3,4) #12 2702 2174 2165 1134
wire n2683; //CHANY (3,4) #13 2663 2084 2059 1134
wire n2684; //CHANY (3,4) #14 2704 2172 2167 1138 890
wire n2685; //CHANY (3,4) #15 2665 2086 2057 1138 890
wire n2686; //CHANY (3,4) #16 2706 2170 2169 894
wire n2687; //CHANY (3,4) #17 2667 2088 2055 894
wire n2688; //CHANY (3,4) #18 2708 2188 2151 1142
wire n2689; //CHANY (3,4) #19 2669 2070 2053 1142
wire n2690; //CHANY (3,5) #0 2270 2251 916
wire n2691; //CHANY (3,5) #1 2671 2172 2151 916
wire n2692; //CHANY (3,5) #2 2272 2253 1164
wire n2693; //CHANY (3,5) #3 2673 2174 2169 1164
wire n2694; //CHANY (3,5) #4 2274 2255 1168 920
wire n2695; //CHANY (3,5) #5 2675 2176 2167 1168 920
wire n2696; //CHANY (3,5) #6 2276 2257 924
wire n2697; //CHANY (3,5) #7 2677 2178 2165 924
wire n2698; //CHANY (3,5) #8 2278 2259 1172
wire n2699; //CHANY (3,5) #9 2679 2180 2163 1172
wire n2700; //CHANY (3,5) #10 2280 2261 916
wire n2701; //CHANY (3,5) #11 2681 2182 2161 916
wire n2702; //CHANY (3,5) #12 2282 2263 1164
wire n2703; //CHANY (3,5) #13 2683 2184 2159 1164
wire n2704; //CHANY (3,5) #14 2284 2265 1168 920
wire n2705; //CHANY (3,5) #15 2685 2186 2157 1168 920
wire n2706; //CHANY (3,5) #16 2286 2267 924
wire n2707; //CHANY (3,5) #17 2687 2188 2155 924
wire n2708; //CHANY (3,5) #18 2288 2269 1172
wire n2709; //CHANY (3,5) #19 2689 2170 2153 1172
wire n2710; //CHANY (4,1) #0 2730 1906 1873 1042
wire n2711; //CHANY (4,1) #1 1790 1771 1042
wire n2712; //CHANY (4,1) #2 2732 1904 1875 1290
wire n2713; //CHANY (4,1) #3 1792 1773 1290
wire n2714; //CHANY (4,1) #4 2734 1902 1877 1294 1046
wire n2715; //CHANY (4,1) #5 1794 1775 1294 1046
wire n2716; //CHANY (4,1) #6 2736 1900 1879 1050
wire n2717; //CHANY (4,1) #7 1796 1777 1050
wire n2718; //CHANY (4,1) #8 2738 1898 1881 1298
wire n2719; //CHANY (4,1) #9 1798 1779 1298
wire n2720; //CHANY (4,1) #10 2740 1896 1883 1042
wire n2721; //CHANY (4,1) #11 1800 1781 1042
wire n2722; //CHANY (4,1) #12 2742 1894 1885 1290
wire n2723; //CHANY (4,1) #13 1802 1783 1290
wire n2724; //CHANY (4,1) #14 2744 1892 1887 1294 1046
wire n2725; //CHANY (4,1) #15 1804 1785 1294 1046
wire n2726; //CHANY (4,1) #16 2746 1890 1889 1050
wire n2727; //CHANY (4,1) #17 1806 1787 1050
wire n2728; //CHANY (4,1) #18 2748 1908 1871 1298
wire n2729; //CHANY (4,1) #19 1808 1789 1298
wire n2730; //CHANY (4,2) #0 2750 2006 1973 1072
wire n2731; //CHANY (4,2) #1 2711 1892 1871 1072
wire n2732; //CHANY (4,2) #2 2752 2004 1975 1320
wire n2733; //CHANY (4,2) #3 2713 1894 1889 1320
wire n2734; //CHANY (4,2) #4 2754 2002 1977 1324 1076
wire n2735; //CHANY (4,2) #5 2715 1896 1887 1324 1076
wire n2736; //CHANY (4,2) #6 2756 2000 1979 1080
wire n2737; //CHANY (4,2) #7 2717 1898 1885 1080
wire n2738; //CHANY (4,2) #8 2758 1998 1981 1328
wire n2739; //CHANY (4,2) #9 2719 1900 1883 1328
wire n2740; //CHANY (4,2) #10 2760 1996 1983 1072
wire n2741; //CHANY (4,2) #11 2721 1902 1881 1072
wire n2742; //CHANY (4,2) #12 2762 1994 1985 1320
wire n2743; //CHANY (4,2) #13 2723 1904 1879 1320
wire n2744; //CHANY (4,2) #14 2764 1992 1987 1324 1076
wire n2745; //CHANY (4,2) #15 2725 1906 1877 1324 1076
wire n2746; //CHANY (4,2) #16 2766 1990 1989 1080
wire n2747; //CHANY (4,2) #17 2727 1908 1875 1080
wire n2748; //CHANY (4,2) #18 2768 2008 1971 1328
wire n2749; //CHANY (4,2) #19 2729 1890 1873 1328
wire n2750; //CHANY (4,3) #0 2770 2106 2073 1102
wire n2751; //CHANY (4,3) #1 2731 1992 1971 1102
wire n2752; //CHANY (4,3) #2 2772 2104 2075 1350
wire n2753; //CHANY (4,3) #3 2733 1994 1989 1350
wire n2754; //CHANY (4,3) #4 2774 2102 2077 1354 1106
wire n2755; //CHANY (4,3) #5 2735 1996 1987 1354 1106
wire n2756; //CHANY (4,3) #6 2776 2100 2079 1110
wire n2757; //CHANY (4,3) #7 2737 1998 1985 1110
wire n2758; //CHANY (4,3) #8 2778 2098 2081 1358
wire n2759; //CHANY (4,3) #9 2739 2000 1983 1358
wire n2760; //CHANY (4,3) #10 2780 2096 2083 1102
wire n2761; //CHANY (4,3) #11 2741 2002 1981 1102
wire n2762; //CHANY (4,3) #12 2782 2094 2085 1350
wire n2763; //CHANY (4,3) #13 2743 2004 1979 1350
wire n2764; //CHANY (4,3) #14 2784 2092 2087 1354 1106
wire n2765; //CHANY (4,3) #15 2745 2006 1977 1354 1106
wire n2766; //CHANY (4,3) #16 2786 2090 2089 1110
wire n2767; //CHANY (4,3) #17 2747 2008 1975 1110
wire n2768; //CHANY (4,3) #18 2788 2108 2071 1358
wire n2769; //CHANY (4,3) #19 2749 1990 1973 1358
wire n2770; //CHANY (4,4) #0 2790 2206 2173 1132
wire n2771; //CHANY (4,4) #1 2751 2092 2071 1132
wire n2772; //CHANY (4,4) #2 2792 2204 2175 1380
wire n2773; //CHANY (4,4) #3 2753 2094 2089 1380
wire n2774; //CHANY (4,4) #4 2794 2202 2177 1384 1136
wire n2775; //CHANY (4,4) #5 2755 2096 2087 1384 1136
wire n2776; //CHANY (4,4) #6 2796 2200 2179 1140
wire n2777; //CHANY (4,4) #7 2757 2098 2085 1140
wire n2778; //CHANY (4,4) #8 2798 2198 2181 1388
wire n2779; //CHANY (4,4) #9 2759 2100 2083 1388
wire n2780; //CHANY (4,4) #10 2800 2196 2183 1132
wire n2781; //CHANY (4,4) #11 2761 2102 2081 1132
wire n2782; //CHANY (4,4) #12 2802 2194 2185 1380
wire n2783; //CHANY (4,4) #13 2763 2104 2079 1380
wire n2784; //CHANY (4,4) #14 2804 2192 2187 1384 1136
wire n2785; //CHANY (4,4) #15 2765 2106 2077 1384 1136
wire n2786; //CHANY (4,4) #16 2806 2190 2189 1140
wire n2787; //CHANY (4,4) #17 2767 2108 2075 1140
wire n2788; //CHANY (4,4) #18 2808 2208 2171 1388
wire n2789; //CHANY (4,4) #19 2769 2090 2073 1388
wire n2790; //CHANY (4,5) #0 2290 2271 1162
wire n2791; //CHANY (4,5) #1 2771 2192 2171 1162
wire n2792; //CHANY (4,5) #2 2292 2273 1410
wire n2793; //CHANY (4,5) #3 2773 2194 2189 1410
wire n2794; //CHANY (4,5) #4 2294 2275 1414 1166
wire n2795; //CHANY (4,5) #5 2775 2196 2187 1414 1166
wire n2796; //CHANY (4,5) #6 2296 2277 1170
wire n2797; //CHANY (4,5) #7 2777 2198 2185 1170
wire n2798; //CHANY (4,5) #8 2298 2279 1418
wire n2799; //CHANY (4,5) #9 2779 2200 2183 1418
wire n2800; //CHANY (4,5) #10 2300 2281 1162
wire n2801; //CHANY (4,5) #11 2781 2202 2181 1162
wire n2802; //CHANY (4,5) #12 2302 2283 1410
wire n2803; //CHANY (4,5) #13 2783 2204 2179 1410
wire n2804; //CHANY (4,5) #14 2304 2285 1414 1166
wire n2805; //CHANY (4,5) #15 2785 2206 2177 1414 1166
wire n2806; //CHANY (4,5) #16 2306 2287 1170
wire n2807; //CHANY (4,5) #17 2787 2208 2175 1170
wire n2808; //CHANY (4,5) #18 2308 2289 1418
wire n2809; //CHANY (4,5) #19 2789 2190 2173 1418
wire n2810; //CHANY (5,1) #0 2830 1891 1494 1288
wire n2811; //CHANY (5,1) #1 1791 1494 1288
wire n2812; //CHANY (5,1) #2 2832 1897 1500 1497
wire n2813; //CHANY (5,1) #3 1809 1500 1497
wire n2814; //CHANY (5,1) #4 2834 1903 1506 1503 1292
wire n2815; //CHANY (5,1) #5 1807 1506 1503 1292
wire n2816; //CHANY (5,1) #6 2836 1909 1509 1296
wire n2817; //CHANY (5,1) #7 1805 1509 1296
wire n2818; //CHANY (5,1) #8 2838 1893 1515 1512
wire n2819; //CHANY (5,1) #9 1803 1515 1512
wire n2820; //CHANY (5,1) #10 2840 1895 1494 1288
wire n2821; //CHANY (5,1) #11 1801 1494 1288
wire n2822; //CHANY (5,1) #12 2842 1899 1500 1497
wire n2823; //CHANY (5,1) #13 1799 1500 1497
wire n2824; //CHANY (5,1) #14 2844 1901 1506 1503 1292
wire n2825; //CHANY (5,1) #15 1797 1506 1503 1292
wire n2826; //CHANY (5,1) #16 2846 1905 1509 1296
wire n2827; //CHANY (5,1) #17 1795 1509 1296
wire n2828; //CHANY (5,1) #18 2848 1907 1515 1512
wire n2829; //CHANY (5,1) #19 1793 1515 1512
wire n2830; //CHANY (5,2) #0 2850 1991 1542 1318
wire n2831; //CHANY (5,2) #1 2811 1891 1542 1318
wire n2832; //CHANY (5,2) #2 2852 1997 1548 1545
wire n2833; //CHANY (5,2) #3 2813 1897 1548 1545
wire n2834; //CHANY (5,2) #4 2854 2003 1554 1551 1322
wire n2835; //CHANY (5,2) #5 2815 1903 1554 1551 1322
wire n2836; //CHANY (5,2) #6 2856 2009 1557 1326
wire n2837; //CHANY (5,2) #7 2817 1909 1557 1326
wire n2838; //CHANY (5,2) #8 2858 1993 1563 1560
wire n2839; //CHANY (5,2) #9 2819 1893 1563 1560
wire n2840; //CHANY (5,2) #10 2860 1995 1542 1318
wire n2841; //CHANY (5,2) #11 2821 1895 1542 1318
wire n2842; //CHANY (5,2) #12 2862 1999 1548 1545
wire n2843; //CHANY (5,2) #13 2823 1899 1548 1545
wire n2844; //CHANY (5,2) #14 2864 2001 1554 1551 1322
wire n2845; //CHANY (5,2) #15 2825 1901 1554 1551 1322
wire n2846; //CHANY (5,2) #16 2866 2005 1557 1326
wire n2847; //CHANY (5,2) #17 2827 1905 1557 1326
wire n2848; //CHANY (5,2) #18 2868 2007 1563 1560
wire n2849; //CHANY (5,2) #19 2829 1907 1563 1560
wire n2850; //CHANY (5,3) #0 2870 2091 1590 1348
wire n2851; //CHANY (5,3) #1 2831 1991 1590 1348
wire n2852; //CHANY (5,3) #2 2872 2097 1596 1593
wire n2853; //CHANY (5,3) #3 2833 1997 1596 1593
wire n2854; //CHANY (5,3) #4 2874 2103 1602 1599 1352
wire n2855; //CHANY (5,3) #5 2835 2003 1602 1599 1352
wire n2856; //CHANY (5,3) #6 2876 2109 1605 1356
wire n2857; //CHANY (5,3) #7 2837 2009 1605 1356
wire n2858; //CHANY (5,3) #8 2878 2093 1611 1608
wire n2859; //CHANY (5,3) #9 2839 1993 1611 1608
wire n2860; //CHANY (5,3) #10 2880 2095 1590 1348
wire n2861; //CHANY (5,3) #11 2841 1995 1590 1348
wire n2862; //CHANY (5,3) #12 2882 2099 1596 1593
wire n2863; //CHANY (5,3) #13 2843 1999 1596 1593
wire n2864; //CHANY (5,3) #14 2884 2101 1602 1599 1352
wire n2865; //CHANY (5,3) #15 2845 2001 1602 1599 1352
wire n2866; //CHANY (5,3) #16 2886 2105 1605 1356
wire n2867; //CHANY (5,3) #17 2847 2005 1605 1356
wire n2868; //CHANY (5,3) #18 2888 2107 1611 1608
wire n2869; //CHANY (5,3) #19 2849 2007 1611 1608
wire n2870; //CHANY (5,4) #0 2890 2191 1638 1378
wire n2871; //CHANY (5,4) #1 2851 2091 1638 1378
wire n2872; //CHANY (5,4) #2 2892 2197 1644 1641
wire n2873; //CHANY (5,4) #3 2853 2097 1644 1641
wire n2874; //CHANY (5,4) #4 2894 2203 1650 1647 1382
wire n2875; //CHANY (5,4) #5 2855 2103 1650 1647 1382
wire n2876; //CHANY (5,4) #6 2896 2209 1653 1386
wire n2877; //CHANY (5,4) #7 2857 2109 1653 1386
wire n2878; //CHANY (5,4) #8 2898 2193 1659 1656
wire n2879; //CHANY (5,4) #9 2859 2093 1659 1656
wire n2880; //CHANY (5,4) #10 2900 2195 1638 1378
wire n2881; //CHANY (5,4) #11 2861 2095 1638 1378
wire n2882; //CHANY (5,4) #12 2902 2199 1644 1641
wire n2883; //CHANY (5,4) #13 2863 2099 1644 1641
wire n2884; //CHANY (5,4) #14 2904 2201 1650 1647 1382
wire n2885; //CHANY (5,4) #15 2865 2101 1650 1647 1382
wire n2886; //CHANY (5,4) #16 2906 2205 1653 1386
wire n2887; //CHANY (5,4) #17 2867 2105 1653 1386
wire n2888; //CHANY (5,4) #18 2908 2207 1659 1656
wire n2889; //CHANY (5,4) #19 2869 2107 1659 1656
wire n2890; //CHANY (5,5) #0 2293 1686 1408
wire n2891; //CHANY (5,5) #1 2871 2191 1686 1408
wire n2892; //CHANY (5,5) #2 2295 1692 1689
wire n2893; //CHANY (5,5) #3 2873 2197 1692 1689
wire n2894; //CHANY (5,5) #4 2297 1698 1695 1412
wire n2895; //CHANY (5,5) #5 2875 2203 1698 1695 1412
wire n2896; //CHANY (5,5) #6 2299 1701 1416
wire n2897; //CHANY (5,5) #7 2877 2209 1701 1416
wire n2898; //CHANY (5,5) #8 2301 1707 1704
wire n2899; //CHANY (5,5) #9 2879 2193 1707 1704
wire n2900; //CHANY (5,5) #10 2303 1686 1408
wire n2901; //CHANY (5,5) #11 2881 2195 1686 1408
wire n2902; //CHANY (5,5) #12 2305 1692 1689
wire n2903; //CHANY (5,5) #13 2883 2199 1692 1689
wire n2904; //CHANY (5,5) #14 2307 1698 1695 1412
wire n2905; //CHANY (5,5) #15 2885 2201 1698 1695 1412
wire n2906; //CHANY (5,5) #16 2309 1701 1416
wire n2907; //CHANY (5,5) #17 2887 2205 1701 1416
wire n2908; //CHANY (5,5) #18 2291 1707 1704
wire n2909; //CHANY (5,5) #19 2889 2207 1707 1704


wire [7777:0] config_chain;
wire [7:0]outpad_0_1;
wire [7:0]inpad_0_1;
io io_0_1 ( .outpad(outpad_0_1), .inpad(inpad_0_1), .io_ext(io_0_1_wire), .config_in(config_chain[7:0]) );

wire [7:0]outpad_0_2;
wire [7:0]inpad_0_2;
io io_0_2 ( .outpad(outpad_0_2), .inpad(inpad_0_2), .io_ext(io_0_2_wire), .config_in(config_chain[15:8]) );

wire [7:0]outpad_0_3;
wire [7:0]inpad_0_3;
io io_0_3 ( .outpad(outpad_0_3), .inpad(inpad_0_3), .io_ext(io_0_3_wire), .config_in(config_chain[23:16]) );

wire [7:0]outpad_0_4;
wire [7:0]inpad_0_4;
io io_0_4 ( .outpad(outpad_0_4), .inpad(inpad_0_4), .io_ext(io_0_4_wire), .config_in(config_chain[31:24]) );

wire [7:0]outpad_0_5;
wire [7:0]inpad_0_5;
io io_0_5 ( .outpad(outpad_0_5), .inpad(inpad_0_5), .io_ext(io_0_5_wire), .config_in(config_chain[39:32]) );

wire [7:0]outpad_1_0;
wire [7:0]inpad_1_0;
io io_1_0 ( .outpad(outpad_1_0), .inpad(inpad_1_0), .io_ext(io_1_0_wire), .config_in(config_chain[47:40]) );

wire [11:0]I_1_1;
wire [1:0]O_1_1;
wire [0:0]clk_1_1;
clb clb_1_1 ( .I(I_1_1), .O(O_1_1), .clk(clk_1_1), .config_in(config_chain[225:48]) );

wire [11:0]I_1_2;
wire [1:0]O_1_2;
wire [0:0]clk_1_2;
clb clb_1_2 ( .I(I_1_2), .O(O_1_2), .clk(clk_1_2), .config_in(config_chain[403:226]) );

wire [11:0]I_1_3;
wire [1:0]O_1_3;
wire [0:0]clk_1_3;
clb clb_1_3 ( .I(I_1_3), .O(O_1_3), .clk(clk_1_3), .config_in(config_chain[581:404]) );

wire [11:0]I_1_4;
wire [1:0]O_1_4;
wire [0:0]clk_1_4;
clb clb_1_4 ( .I(I_1_4), .O(O_1_4), .clk(clk_1_4), .config_in(config_chain[759:582]) );

wire [11:0]I_1_5;
wire [1:0]O_1_5;
wire [0:0]clk_1_5;
clb clb_1_5 ( .I(I_1_5), .O(O_1_5), .clk(clk_1_5), .config_in(config_chain[937:760]) );

wire [7:0]outpad_1_6;
wire [7:0]inpad_1_6;
io io_1_6 ( .outpad(outpad_1_6), .inpad(inpad_1_6), .io_ext(io_1_6_wire), .config_in(config_chain[945:938]) );

wire [7:0]outpad_2_0;
wire [7:0]inpad_2_0;
io io_2_0 ( .outpad(outpad_2_0), .inpad(inpad_2_0), .io_ext(io_2_0_wire), .config_in(config_chain[953:946]) );

wire [11:0]I_2_1;
wire [1:0]O_2_1;
wire [0:0]clk_2_1;
clb clb_2_1 ( .I(I_2_1), .O(O_2_1), .clk(clk_2_1), .config_in(config_chain[1131:954]) );

wire [11:0]I_2_2;
wire [1:0]O_2_2;
wire [0:0]clk_2_2;
clb clb_2_2 ( .I(I_2_2), .O(O_2_2), .clk(clk_2_2), .config_in(config_chain[1309:1132]) );

wire [11:0]I_2_3;
wire [1:0]O_2_3;
wire [0:0]clk_2_3;
clb clb_2_3 ( .I(I_2_3), .O(O_2_3), .clk(clk_2_3), .config_in(config_chain[1487:1310]) );

wire [11:0]I_2_4;
wire [1:0]O_2_4;
wire [0:0]clk_2_4;
clb clb_2_4 ( .I(I_2_4), .O(O_2_4), .clk(clk_2_4), .config_in(config_chain[1665:1488]) );

wire [11:0]I_2_5;
wire [1:0]O_2_5;
wire [0:0]clk_2_5;
clb clb_2_5 ( .I(I_2_5), .O(O_2_5), .clk(clk_2_5), .config_in(config_chain[1843:1666]) );

wire [7:0]outpad_2_6;
wire [7:0]inpad_2_6;
io io_2_6 ( .outpad(outpad_2_6), .inpad(inpad_2_6), .io_ext(io_2_6_wire), .config_in(config_chain[1851:1844]) );

wire [7:0]outpad_3_0;
wire [7:0]inpad_3_0;
io io_3_0 ( .outpad(outpad_3_0), .inpad(inpad_3_0), .io_ext(io_3_0_wire), .config_in(config_chain[1859:1852]) );

wire [11:0]I_3_1;
wire [1:0]O_3_1;
wire [0:0]clk_3_1;
clb clb_3_1 ( .I(I_3_1), .O(O_3_1), .clk(clk_3_1), .config_in(config_chain[2037:1860]) );

wire [11:0]I_3_2;
wire [1:0]O_3_2;
wire [0:0]clk_3_2;
clb clb_3_2 ( .I(I_3_2), .O(O_3_2), .clk(clk_3_2), .config_in(config_chain[2215:2038]) );

wire [11:0]I_3_3;
wire [1:0]O_3_3;
wire [0:0]clk_3_3;
clb clb_3_3 ( .I(I_3_3), .O(O_3_3), .clk(clk_3_3), .config_in(config_chain[2393:2216]) );

wire [11:0]I_3_4;
wire [1:0]O_3_4;
wire [0:0]clk_3_4;
clb clb_3_4 ( .I(I_3_4), .O(O_3_4), .clk(clk_3_4), .config_in(config_chain[2571:2394]) );

wire [11:0]I_3_5;
wire [1:0]O_3_5;
wire [0:0]clk_3_5;
clb clb_3_5 ( .I(I_3_5), .O(O_3_5), .clk(clk_3_5), .config_in(config_chain[2749:2572]) );

wire [7:0]outpad_3_6;
wire [7:0]inpad_3_6;
io io_3_6 ( .outpad(outpad_3_6), .inpad(inpad_3_6), .io_ext(io_3_6_wire), .config_in(config_chain[2757:2750]) );

wire [7:0]outpad_4_0;
wire [7:0]inpad_4_0;
io io_4_0 ( .outpad(outpad_4_0), .inpad(inpad_4_0), .io_ext(io_4_0_wire), .config_in(config_chain[2765:2758]) );

wire [11:0]I_4_1;
wire [1:0]O_4_1;
wire [0:0]clk_4_1;
clb clb_4_1 ( .I(I_4_1), .O(O_4_1), .clk(clk_4_1), .config_in(config_chain[2943:2766]) );

wire [11:0]I_4_2;
wire [1:0]O_4_2;
wire [0:0]clk_4_2;
clb clb_4_2 ( .I(I_4_2), .O(O_4_2), .clk(clk_4_2), .config_in(config_chain[3121:2944]) );

wire [11:0]I_4_3;
wire [1:0]O_4_3;
wire [0:0]clk_4_3;
clb clb_4_3 ( .I(I_4_3), .O(O_4_3), .clk(clk_4_3), .config_in(config_chain[3299:3122]) );

wire [11:0]I_4_4;
wire [1:0]O_4_4;
wire [0:0]clk_4_4;
clb clb_4_4 ( .I(I_4_4), .O(O_4_4), .clk(clk_4_4), .config_in(config_chain[3477:3300]) );

wire [11:0]I_4_5;
wire [1:0]O_4_5;
wire [0:0]clk_4_5;
clb clb_4_5 ( .I(I_4_5), .O(O_4_5), .clk(clk_4_5), .config_in(config_chain[3655:3478]) );

wire [7:0]outpad_4_6;
wire [7:0]inpad_4_6;
io io_4_6 ( .outpad(outpad_4_6), .inpad(inpad_4_6), .io_ext(io_4_6_wire), .config_in(config_chain[3663:3656]) );

wire [7:0]outpad_5_0;
wire [7:0]inpad_5_0;
io io_5_0 ( .outpad(outpad_5_0), .inpad(inpad_5_0), .io_ext(io_5_0_wire), .config_in(config_chain[3671:3664]) );

wire [11:0]I_5_1;
wire [1:0]O_5_1;
wire [0:0]clk_5_1;
clb clb_5_1 ( .I(I_5_1), .O(O_5_1), .clk(clk_5_1), .config_in(config_chain[3849:3672]) );

wire [11:0]I_5_2;
wire [1:0]O_5_2;
wire [0:0]clk_5_2;
clb clb_5_2 ( .I(I_5_2), .O(O_5_2), .clk(clk_5_2), .config_in(config_chain[4027:3850]) );

wire [11:0]I_5_3;
wire [1:0]O_5_3;
wire [0:0]clk_5_3;
clb clb_5_3 ( .I(I_5_3), .O(O_5_3), .clk(clk_5_3), .config_in(config_chain[4205:4028]) );

wire [11:0]I_5_4;
wire [1:0]O_5_4;
wire [0:0]clk_5_4;
clb clb_5_4 ( .I(I_5_4), .O(O_5_4), .clk(clk_5_4), .config_in(config_chain[4383:4206]) );

wire [11:0]I_5_5;
wire [1:0]O_5_5;
wire [0:0]clk_5_5;
clb clb_5_5 ( .I(I_5_5), .O(O_5_5), .clk(clk_5_5), .config_in(config_chain[4561:4384]) );

wire [7:0]outpad_5_6;
wire [7:0]inpad_5_6;
io io_5_6 ( .outpad(outpad_5_6), .inpad(inpad_5_6), .io_ext(io_5_6_wire), .config_in(config_chain[4569:4562]) );

wire [7:0]outpad_6_1;
wire [7:0]inpad_6_1;
io io_6_1 ( .outpad(outpad_6_1), .inpad(inpad_6_1), .io_ext(io_6_1_wire), .config_in(config_chain[4577:4570]) );

wire [7:0]outpad_6_2;
wire [7:0]inpad_6_2;
io io_6_2 ( .outpad(outpad_6_2), .inpad(inpad_6_2), .io_ext(io_6_2_wire), .config_in(config_chain[4585:4578]) );

wire [7:0]outpad_6_3;
wire [7:0]inpad_6_3;
io io_6_3 ( .outpad(outpad_6_3), .inpad(inpad_6_3), .io_ext(io_6_3_wire), .config_in(config_chain[4593:4586]) );

wire [7:0]outpad_6_4;
wire [7:0]inpad_6_4;
io io_6_4 ( .outpad(outpad_6_4), .inpad(inpad_6_4), .io_ext(io_6_4_wire), .config_in(config_chain[4601:4594]) );

wire [7:0]outpad_6_5;
wire [7:0]inpad_6_5;
io io_6_5 ( .outpad(outpad_6_5), .inpad(inpad_6_5), .io_ext(io_6_5_wire), .config_in(config_chain[4609:4602]) );

assign outpad_0_1 = {n45, n42, n39, n36, n33, n30, n27, n24};
assign {n46, n43, n40, n37, n34, n31, n28, n25} = inpad_0_1;
assign outpad_0_2 = {n93, n90, n87, n84, n81, n78, n75, n72};
assign {n94, n91, n88, n85, n82, n79, n76, n73} = inpad_0_2;
assign outpad_0_3 = {n141, n138, n135, n132, n129, n126, n123, n120};
assign {n142, n139, n136, n133, n130, n127, n124, n121} = inpad_0_3;
assign outpad_0_4 = {n189, n186, n183, n180, n177, n174, n171, n168};
assign {n190, n187, n184, n181, n178, n175, n172, n169} = inpad_0_4;
assign outpad_0_5 = {n237, n234, n231, n228, n225, n222, n219, n216};
assign {n238, n235, n232, n229, n226, n223, n220, n217} = inpad_0_5;
assign outpad_1_0 = {n285, n282, n279, n276, n273, n270, n267, n264};
assign {n286, n283, n280, n277, n274, n271, n268, n265} = inpad_1_0;
assign clk_1_1 = {clk};
assign I_1_1 = {n314, n313, n312, n311, n310, n309, n308, n307, n306, n305, n304, n303};
assign {n316, n315} = O_1_1;
assign clk_1_2 = {clk};
assign I_1_2 = {n344, n343, n342, n341, n340, n339, n338, n337, n336, n335, n334, n333};
assign {n346, n345} = O_1_2;
assign clk_1_3 = {clk};
assign I_1_3 = {n374, n373, n372, n371, n370, n369, n368, n367, n366, n365, n364, n363};
assign {n376, n375} = O_1_3;
assign clk_1_4 = {clk};
assign I_1_4 = {n404, n403, n402, n401, n400, n399, n398, n397, n396, n395, n394, n393};
assign {n406, n405} = O_1_4;
assign clk_1_5 = {clk};
assign I_1_5 = {n434, n433, n432, n431, n430, n429, n428, n427, n426, n425, n424, n423};
assign {n436, n435} = O_1_5;
assign outpad_1_6 = {n483, n480, n477, n474, n471, n468, n465, n462};
assign {n484, n481, n478, n475, n472, n469, n466, n463} = inpad_1_6;
assign outpad_2_0 = {n531, n528, n525, n522, n519, n516, n513, n510};
assign {n532, n529, n526, n523, n520, n517, n514, n511} = inpad_2_0;
assign clk_2_1 = {clk};
assign I_2_1 = {n560, n559, n558, n557, n556, n555, n554, n553, n552, n551, n550, n549};
assign {n562, n561} = O_2_1;
assign clk_2_2 = {clk};
assign I_2_2 = {n590, n589, n588, n587, n586, n585, n584, n583, n582, n581, n580, n579};
assign {n592, n591} = O_2_2;
assign clk_2_3 = {clk};
assign I_2_3 = {n620, n619, n618, n617, n616, n615, n614, n613, n612, n611, n610, n609};
assign {n622, n621} = O_2_3;
assign clk_2_4 = {clk};
assign I_2_4 = {n650, n649, n648, n647, n646, n645, n644, n643, n642, n641, n640, n639};
assign {n652, n651} = O_2_4;
assign clk_2_5 = {clk};
assign I_2_5 = {n680, n679, n678, n677, n676, n675, n674, n673, n672, n671, n670, n669};
assign {n682, n681} = O_2_5;
assign outpad_2_6 = {n729, n726, n723, n720, n717, n714, n711, n708};
assign {n730, n727, n724, n721, n718, n715, n712, n709} = inpad_2_6;
assign outpad_3_0 = {n777, n774, n771, n768, n765, n762, n759, n756};
assign {n778, n775, n772, n769, n766, n763, n760, n757} = inpad_3_0;
assign clk_3_1 = {clk};
assign I_3_1 = {n806, n805, n804, n803, n802, n801, n800, n799, n798, n797, n796, n795};
assign {n808, n807} = O_3_1;
assign clk_3_2 = {clk};
assign I_3_2 = {n836, n835, n834, n833, n832, n831, n830, n829, n828, n827, n826, n825};
assign {n838, n837} = O_3_2;
assign clk_3_3 = {clk};
assign I_3_3 = {n866, n865, n864, n863, n862, n861, n860, n859, n858, n857, n856, n855};
assign {n868, n867} = O_3_3;
assign clk_3_4 = {clk};
assign I_3_4 = {n896, n895, n894, n893, n892, n891, n890, n889, n888, n887, n886, n885};
assign {n898, n897} = O_3_4;
assign clk_3_5 = {clk};
assign I_3_5 = {n926, n925, n924, n923, n922, n921, n920, n919, n918, n917, n916, n915};
assign {n928, n927} = O_3_5;
assign outpad_3_6 = {n975, n972, n969, n966, n963, n960, n957, n954};
assign {n976, n973, n970, n967, n964, n961, n958, n955} = inpad_3_6;
assign outpad_4_0 = {n1023, n1020, n1017, n1014, n1011, n1008, n1005, n1002};
assign {n1024, n1021, n1018, n1015, n1012, n1009, n1006, n1003} = inpad_4_0;
assign clk_4_1 = {clk};
assign I_4_1 = {n1052, n1051, n1050, n1049, n1048, n1047, n1046, n1045, n1044, n1043, n1042, n1041};
assign {n1054, n1053} = O_4_1;
assign clk_4_2 = {clk};
assign I_4_2 = {n1082, n1081, n1080, n1079, n1078, n1077, n1076, n1075, n1074, n1073, n1072, n1071};
assign {n1084, n1083} = O_4_2;
assign clk_4_3 = {clk};
assign I_4_3 = {n1112, n1111, n1110, n1109, n1108, n1107, n1106, n1105, n1104, n1103, n1102, n1101};
assign {n1114, n1113} = O_4_3;
assign clk_4_4 = {clk};
assign I_4_4 = {n1142, n1141, n1140, n1139, n1138, n1137, n1136, n1135, n1134, n1133, n1132, n1131};
assign {n1144, n1143} = O_4_4;
assign clk_4_5 = {clk};
assign I_4_5 = {n1172, n1171, n1170, n1169, n1168, n1167, n1166, n1165, n1164, n1163, n1162, n1161};
assign {n1174, n1173} = O_4_5;
assign outpad_4_6 = {n1221, n1218, n1215, n1212, n1209, n1206, n1203, n1200};
assign {n1222, n1219, n1216, n1213, n1210, n1207, n1204, n1201} = inpad_4_6;
assign outpad_5_0 = {n1269, n1266, n1263, n1260, n1257, n1254, n1251, n1248};
assign {n1270, n1267, n1264, n1261, n1258, n1255, n1252, n1249} = inpad_5_0;
assign clk_5_1 = {clk};
assign I_5_1 = {n1298, n1297, n1296, n1295, n1294, n1293, n1292, n1291, n1290, n1289, n1288, n1287};
assign {n1300, n1299} = O_5_1;
assign clk_5_2 = {clk};
assign I_5_2 = {n1328, n1327, n1326, n1325, n1324, n1323, n1322, n1321, n1320, n1319, n1318, n1317};
assign {n1330, n1329} = O_5_2;
assign clk_5_3 = {clk};
assign I_5_3 = {n1358, n1357, n1356, n1355, n1354, n1353, n1352, n1351, n1350, n1349, n1348, n1347};
assign {n1360, n1359} = O_5_3;
assign clk_5_4 = {clk};
assign I_5_4 = {n1388, n1387, n1386, n1385, n1384, n1383, n1382, n1381, n1380, n1379, n1378, n1377};
assign {n1390, n1389} = O_5_4;
assign clk_5_5 = {clk};
assign I_5_5 = {n1418, n1417, n1416, n1415, n1414, n1413, n1412, n1411, n1410, n1409, n1408, n1407};
assign {n1420, n1419} = O_5_5;
assign outpad_5_6 = {n1467, n1464, n1461, n1458, n1455, n1452, n1449, n1446};
assign {n1468, n1465, n1462, n1459, n1456, n1453, n1450, n1447} = inpad_5_6;
assign outpad_6_1 = {n1515, n1512, n1509, n1506, n1503, n1500, n1497, n1494};
assign {n1516, n1513, n1510, n1507, n1504, n1501, n1498, n1495} = inpad_6_1;
assign outpad_6_2 = {n1563, n1560, n1557, n1554, n1551, n1548, n1545, n1542};
assign {n1564, n1561, n1558, n1555, n1552, n1549, n1546, n1543} = inpad_6_2;
assign outpad_6_3 = {n1611, n1608, n1605, n1602, n1599, n1596, n1593, n1590};
assign {n1612, n1609, n1606, n1603, n1600, n1597, n1594, n1591} = inpad_6_3;
assign outpad_6_4 = {n1659, n1656, n1653, n1650, n1647, n1644, n1641, n1638};
assign {n1660, n1657, n1654, n1651, n1648, n1645, n1642, n1639} = inpad_6_4;
assign outpad_6_5 = {n1707, n1704, n1701, n1698, n1695, n1692, n1689, n1686};
assign {n1708, n1705, n1702, n1699, n1696, n1693, n1690, n1687} = inpad_6_5;

mux4 mux_0 (.in({n2321, n2320, n2311, n2310}), .out(n24), .config_in(config_chain[4611:4610])); 
mux4 mux_1 (.in({n2321, n2320, n2311, n2310}), .out(n27), .config_in(config_chain[4613:4612])); 
mux4 mux_2 (.in({n2323, n2322, n2313, n2312}), .out(n30), .config_in(config_chain[4615:4614])); 
mux4 mux_3 (.in({n2325, n2324, n2315, n2314}), .out(n33), .config_in(config_chain[4617:4616])); 
mux4 mux_4 (.in({n2325, n2324, n2315, n2314}), .out(n36), .config_in(config_chain[4619:4618])); 
mux4 mux_5 (.in({n2327, n2326, n2317, n2316}), .out(n39), .config_in(config_chain[4621:4620])); 
mux4 mux_6 (.in({n2327, n2326, n2317, n2316}), .out(n42), .config_in(config_chain[4623:4622])); 
mux4 mux_7 (.in({n2329, n2328, n2319, n2318}), .out(n45), .config_in(config_chain[4625:4624])); 
mux4 mux_8 (.in({n2341, n2340, n2331, n2330}), .out(n72), .config_in(config_chain[4627:4626])); 
mux4 mux_9 (.in({n2341, n2340, n2331, n2330}), .out(n75), .config_in(config_chain[4629:4628])); 
mux4 mux_10 (.in({n2343, n2342, n2333, n2332}), .out(n78), .config_in(config_chain[4631:4630])); 
mux4 mux_11 (.in({n2345, n2344, n2335, n2334}), .out(n81), .config_in(config_chain[4633:4632])); 
mux4 mux_12 (.in({n2345, n2344, n2335, n2334}), .out(n84), .config_in(config_chain[4635:4634])); 
mux4 mux_13 (.in({n2347, n2346, n2337, n2336}), .out(n87), .config_in(config_chain[4637:4636])); 
mux4 mux_14 (.in({n2347, n2346, n2337, n2336}), .out(n90), .config_in(config_chain[4639:4638])); 
mux4 mux_15 (.in({n2349, n2348, n2339, n2338}), .out(n93), .config_in(config_chain[4641:4640])); 
mux4 mux_16 (.in({n2361, n2360, n2351, n2350}), .out(n120), .config_in(config_chain[4643:4642])); 
mux4 mux_17 (.in({n2361, n2360, n2351, n2350}), .out(n123), .config_in(config_chain[4645:4644])); 
mux4 mux_18 (.in({n2363, n2362, n2353, n2352}), .out(n126), .config_in(config_chain[4647:4646])); 
mux4 mux_19 (.in({n2365, n2364, n2355, n2354}), .out(n129), .config_in(config_chain[4649:4648])); 
mux4 mux_20 (.in({n2365, n2364, n2355, n2354}), .out(n132), .config_in(config_chain[4651:4650])); 
mux4 mux_21 (.in({n2367, n2366, n2357, n2356}), .out(n135), .config_in(config_chain[4653:4652])); 
mux4 mux_22 (.in({n2367, n2366, n2357, n2356}), .out(n138), .config_in(config_chain[4655:4654])); 
mux4 mux_23 (.in({n2369, n2368, n2359, n2358}), .out(n141), .config_in(config_chain[4657:4656])); 
mux4 mux_24 (.in({n2381, n2380, n2371, n2370}), .out(n168), .config_in(config_chain[4659:4658])); 
mux4 mux_25 (.in({n2381, n2380, n2371, n2370}), .out(n171), .config_in(config_chain[4661:4660])); 
mux4 mux_26 (.in({n2383, n2382, n2373, n2372}), .out(n174), .config_in(config_chain[4663:4662])); 
mux4 mux_27 (.in({n2385, n2384, n2375, n2374}), .out(n177), .config_in(config_chain[4665:4664])); 
mux4 mux_28 (.in({n2385, n2384, n2375, n2374}), .out(n180), .config_in(config_chain[4667:4666])); 
mux4 mux_29 (.in({n2387, n2386, n2377, n2376}), .out(n183), .config_in(config_chain[4669:4668])); 
mux4 mux_30 (.in({n2387, n2386, n2377, n2376}), .out(n186), .config_in(config_chain[4671:4670])); 
mux4 mux_31 (.in({n2389, n2388, n2379, n2378}), .out(n189), .config_in(config_chain[4673:4672])); 
mux4 mux_32 (.in({n2401, n2400, n2391, n2390}), .out(n216), .config_in(config_chain[4675:4674])); 
mux4 mux_33 (.in({n2401, n2400, n2391, n2390}), .out(n219), .config_in(config_chain[4677:4676])); 
mux4 mux_34 (.in({n2403, n2402, n2393, n2392}), .out(n222), .config_in(config_chain[4679:4678])); 
mux4 mux_35 (.in({n2405, n2404, n2395, n2394}), .out(n225), .config_in(config_chain[4681:4680])); 
mux4 mux_36 (.in({n2405, n2404, n2395, n2394}), .out(n228), .config_in(config_chain[4683:4682])); 
mux4 mux_37 (.in({n2407, n2406, n2397, n2396}), .out(n231), .config_in(config_chain[4685:4684])); 
mux4 mux_38 (.in({n2407, n2406, n2397, n2396}), .out(n234), .config_in(config_chain[4687:4686])); 
mux4 mux_39 (.in({n2409, n2408, n2399, n2398}), .out(n237), .config_in(config_chain[4689:4688])); 
mux4 mux_40 (.in({n1721, n1720, n1711, n1710}), .out(n264), .config_in(config_chain[4691:4690])); 
mux4 mux_41 (.in({n1721, n1720, n1711, n1710}), .out(n267), .config_in(config_chain[4693:4692])); 
mux4 mux_42 (.in({n1723, n1722, n1713, n1712}), .out(n270), .config_in(config_chain[4695:4694])); 
mux4 mux_43 (.in({n1723, n1722, n1713, n1712}), .out(n273), .config_in(config_chain[4697:4696])); 
mux4 mux_44 (.in({n1725, n1724, n1715, n1714}), .out(n276), .config_in(config_chain[4699:4698])); 
mux4 mux_45 (.in({n1727, n1726, n1717, n1716}), .out(n279), .config_in(config_chain[4701:4700])); 
mux4 mux_46 (.in({n1727, n1726, n1717, n1716}), .out(n282), .config_in(config_chain[4703:4702])); 
mux4 mux_47 (.in({n1729, n1728, n1719, n1718}), .out(n285), .config_in(config_chain[4705:4704])); 
mux4 mux_48 (.in({n1821, n1820, n1811, n1810}), .out(n303), .config_in(config_chain[4707:4706])); 
mux4 mux_49 (.in({n2421, n2420, n2411, n2410}), .out(n304), .config_in(config_chain[4709:4708])); 
mux4 mux_50 (.in({n1721, n1720, n1711, n1710}), .out(n305), .config_in(config_chain[4711:4710])); 
mux4 mux_51 (.in({n2323, n2322, n2313, n2312}), .out(n306), .config_in(config_chain[4713:4712])); 
mux4 mux_52 (.in({n1823, n1822, n1813, n1812}), .out(n307), .config_in(config_chain[4715:4714])); 
mux4 mux_53 (.in({n2425, n2424, n2415, n2414}), .out(n308), .config_in(config_chain[4717:4716])); 
mux4 mux_54 (.in({n1725, n1724, n1715, n1714}), .out(n309), .config_in(config_chain[4719:4718])); 
mux4 mux_55 (.in({n2325, n2324, n2315, n2314}), .out(n310), .config_in(config_chain[4721:4720])); 
mux4 mux_56 (.in({n1827, n1826, n1817, n1816}), .out(n311), .config_in(config_chain[4723:4722])); 
mux4 mux_57 (.in({n2427, n2426, n2417, n2416}), .out(n312), .config_in(config_chain[4725:4724])); 
mux4 mux_58 (.in({n1729, n1728, n1719, n1718}), .out(n313), .config_in(config_chain[4727:4726])); 
mux4 mux_59 (.in({n2329, n2328, n2319, n2318}), .out(n314), .config_in(config_chain[4729:4728])); 
mux4 mux_60 (.in({n1921, n1920, n1911, n1910}), .out(n333), .config_in(config_chain[4731:4730])); 
mux4 mux_61 (.in({n2441, n2440, n2431, n2430}), .out(n334), .config_in(config_chain[4733:4732])); 
mux4 mux_62 (.in({n1821, n1820, n1811, n1810}), .out(n335), .config_in(config_chain[4735:4734])); 
mux4 mux_63 (.in({n2343, n2342, n2333, n2332}), .out(n336), .config_in(config_chain[4737:4736])); 
mux4 mux_64 (.in({n1923, n1922, n1913, n1912}), .out(n337), .config_in(config_chain[4739:4738])); 
mux4 mux_65 (.in({n2445, n2444, n2435, n2434}), .out(n338), .config_in(config_chain[4741:4740])); 
mux4 mux_66 (.in({n1825, n1824, n1815, n1814}), .out(n339), .config_in(config_chain[4743:4742])); 
mux4 mux_67 (.in({n2345, n2344, n2335, n2334}), .out(n340), .config_in(config_chain[4745:4744])); 
mux4 mux_68 (.in({n1927, n1926, n1917, n1916}), .out(n341), .config_in(config_chain[4747:4746])); 
mux4 mux_69 (.in({n2447, n2446, n2437, n2436}), .out(n342), .config_in(config_chain[4749:4748])); 
mux4 mux_70 (.in({n1829, n1828, n1819, n1818}), .out(n343), .config_in(config_chain[4751:4750])); 
mux4 mux_71 (.in({n2349, n2348, n2339, n2338}), .out(n344), .config_in(config_chain[4753:4752])); 
mux4 mux_72 (.in({n2021, n2020, n2011, n2010}), .out(n363), .config_in(config_chain[4755:4754])); 
mux4 mux_73 (.in({n2461, n2460, n2451, n2450}), .out(n364), .config_in(config_chain[4757:4756])); 
mux4 mux_74 (.in({n1921, n1920, n1911, n1910}), .out(n365), .config_in(config_chain[4759:4758])); 
mux4 mux_75 (.in({n2363, n2362, n2353, n2352}), .out(n366), .config_in(config_chain[4761:4760])); 
mux4 mux_76 (.in({n2023, n2022, n2013, n2012}), .out(n367), .config_in(config_chain[4763:4762])); 
mux4 mux_77 (.in({n2465, n2464, n2455, n2454}), .out(n368), .config_in(config_chain[4765:4764])); 
mux4 mux_78 (.in({n1925, n1924, n1915, n1914}), .out(n369), .config_in(config_chain[4767:4766])); 
mux4 mux_79 (.in({n2365, n2364, n2355, n2354}), .out(n370), .config_in(config_chain[4769:4768])); 
mux4 mux_80 (.in({n2027, n2026, n2017, n2016}), .out(n371), .config_in(config_chain[4771:4770])); 
mux4 mux_81 (.in({n2467, n2466, n2457, n2456}), .out(n372), .config_in(config_chain[4773:4772])); 
mux4 mux_82 (.in({n1929, n1928, n1919, n1918}), .out(n373), .config_in(config_chain[4775:4774])); 
mux4 mux_83 (.in({n2369, n2368, n2359, n2358}), .out(n374), .config_in(config_chain[4777:4776])); 
mux4 mux_84 (.in({n2121, n2120, n2111, n2110}), .out(n393), .config_in(config_chain[4779:4778])); 
mux4 mux_85 (.in({n2481, n2480, n2471, n2470}), .out(n394), .config_in(config_chain[4781:4780])); 
mux4 mux_86 (.in({n2021, n2020, n2011, n2010}), .out(n395), .config_in(config_chain[4783:4782])); 
mux4 mux_87 (.in({n2383, n2382, n2373, n2372}), .out(n396), .config_in(config_chain[4785:4784])); 
mux4 mux_88 (.in({n2123, n2122, n2113, n2112}), .out(n397), .config_in(config_chain[4787:4786])); 
mux4 mux_89 (.in({n2485, n2484, n2475, n2474}), .out(n398), .config_in(config_chain[4789:4788])); 
mux4 mux_90 (.in({n2025, n2024, n2015, n2014}), .out(n399), .config_in(config_chain[4791:4790])); 
mux4 mux_91 (.in({n2385, n2384, n2375, n2374}), .out(n400), .config_in(config_chain[4793:4792])); 
mux4 mux_92 (.in({n2127, n2126, n2117, n2116}), .out(n401), .config_in(config_chain[4795:4794])); 
mux4 mux_93 (.in({n2487, n2486, n2477, n2476}), .out(n402), .config_in(config_chain[4797:4796])); 
mux4 mux_94 (.in({n2029, n2028, n2019, n2018}), .out(n403), .config_in(config_chain[4799:4798])); 
mux4 mux_95 (.in({n2389, n2388, n2379, n2378}), .out(n404), .config_in(config_chain[4801:4800])); 
mux4 mux_96 (.in({n2221, n2220, n2211, n2210}), .out(n423), .config_in(config_chain[4803:4802])); 
mux4 mux_97 (.in({n2501, n2500, n2491, n2490}), .out(n424), .config_in(config_chain[4805:4804])); 
mux4 mux_98 (.in({n2121, n2120, n2111, n2110}), .out(n425), .config_in(config_chain[4807:4806])); 
mux4 mux_99 (.in({n2403, n2402, n2393, n2392}), .out(n426), .config_in(config_chain[4809:4808])); 
mux4 mux_100 (.in({n2223, n2222, n2213, n2212}), .out(n427), .config_in(config_chain[4811:4810])); 
mux4 mux_101 (.in({n2505, n2504, n2495, n2494}), .out(n428), .config_in(config_chain[4813:4812])); 
mux4 mux_102 (.in({n2125, n2124, n2115, n2114}), .out(n429), .config_in(config_chain[4815:4814])); 
mux4 mux_103 (.in({n2405, n2404, n2395, n2394}), .out(n430), .config_in(config_chain[4817:4816])); 
mux4 mux_104 (.in({n2227, n2226, n2217, n2216}), .out(n431), .config_in(config_chain[4819:4818])); 
mux4 mux_105 (.in({n2507, n2506, n2497, n2496}), .out(n432), .config_in(config_chain[4821:4820])); 
mux4 mux_106 (.in({n2129, n2128, n2119, n2118}), .out(n433), .config_in(config_chain[4823:4822])); 
mux4 mux_107 (.in({n2409, n2408, n2399, n2398}), .out(n434), .config_in(config_chain[4825:4824])); 
mux4 mux_108 (.in({n2221, n2220, n2211, n2210}), .out(n462), .config_in(config_chain[4827:4826])); 
mux4 mux_109 (.in({n2221, n2220, n2211, n2210}), .out(n465), .config_in(config_chain[4829:4828])); 
mux4 mux_110 (.in({n2223, n2222, n2213, n2212}), .out(n468), .config_in(config_chain[4831:4830])); 
mux4 mux_111 (.in({n2225, n2224, n2215, n2214}), .out(n471), .config_in(config_chain[4833:4832])); 
mux4 mux_112 (.in({n2225, n2224, n2215, n2214}), .out(n474), .config_in(config_chain[4835:4834])); 
mux4 mux_113 (.in({n2227, n2226, n2217, n2216}), .out(n477), .config_in(config_chain[4837:4836])); 
mux4 mux_114 (.in({n2229, n2228, n2219, n2218}), .out(n480), .config_in(config_chain[4839:4838])); 
mux4 mux_115 (.in({n2229, n2228, n2219, n2218}), .out(n483), .config_in(config_chain[4841:4840])); 
mux4 mux_116 (.in({n1741, n1740, n1731, n1730}), .out(n510), .config_in(config_chain[4843:4842])); 
mux4 mux_117 (.in({n1741, n1740, n1731, n1730}), .out(n513), .config_in(config_chain[4845:4844])); 
mux4 mux_118 (.in({n1743, n1742, n1733, n1732}), .out(n516), .config_in(config_chain[4847:4846])); 
mux4 mux_119 (.in({n1743, n1742, n1733, n1732}), .out(n519), .config_in(config_chain[4849:4848])); 
mux4 mux_120 (.in({n1745, n1744, n1735, n1734}), .out(n522), .config_in(config_chain[4851:4850])); 
mux4 mux_121 (.in({n1747, n1746, n1737, n1736}), .out(n525), .config_in(config_chain[4853:4852])); 
mux4 mux_122 (.in({n1747, n1746, n1737, n1736}), .out(n528), .config_in(config_chain[4855:4854])); 
mux4 mux_123 (.in({n1749, n1748, n1739, n1738}), .out(n531), .config_in(config_chain[4857:4856])); 
mux4 mux_124 (.in({n1841, n1840, n1831, n1830}), .out(n549), .config_in(config_chain[4859:4858])); 
mux4 mux_125 (.in({n2521, n2520, n2511, n2510}), .out(n550), .config_in(config_chain[4861:4860])); 
mux4 mux_126 (.in({n1741, n1740, n1731, n1730}), .out(n551), .config_in(config_chain[4863:4862])); 
mux4 mux_127 (.in({n2423, n2422, n2413, n2412}), .out(n552), .config_in(config_chain[4865:4864])); 
mux4 mux_128 (.in({n1843, n1842, n1833, n1832}), .out(n553), .config_in(config_chain[4867:4866])); 
mux4 mux_129 (.in({n2525, n2524, n2515, n2514}), .out(n554), .config_in(config_chain[4869:4868])); 
mux4 mux_130 (.in({n1745, n1744, n1735, n1734}), .out(n555), .config_in(config_chain[4871:4870])); 
mux4 mux_131 (.in({n2425, n2424, n2415, n2414}), .out(n556), .config_in(config_chain[4873:4872])); 
mux4 mux_132 (.in({n1847, n1846, n1837, n1836}), .out(n557), .config_in(config_chain[4875:4874])); 
mux4 mux_133 (.in({n2527, n2526, n2517, n2516}), .out(n558), .config_in(config_chain[4877:4876])); 
mux4 mux_134 (.in({n1749, n1748, n1739, n1738}), .out(n559), .config_in(config_chain[4879:4878])); 
mux4 mux_135 (.in({n2429, n2428, n2419, n2418}), .out(n560), .config_in(config_chain[4881:4880])); 
mux4 mux_136 (.in({n1941, n1940, n1931, n1930}), .out(n579), .config_in(config_chain[4883:4882])); 
mux4 mux_137 (.in({n2541, n2540, n2531, n2530}), .out(n580), .config_in(config_chain[4885:4884])); 
mux4 mux_138 (.in({n1841, n1840, n1831, n1830}), .out(n581), .config_in(config_chain[4887:4886])); 
mux4 mux_139 (.in({n2443, n2442, n2433, n2432}), .out(n582), .config_in(config_chain[4889:4888])); 
mux4 mux_140 (.in({n1943, n1942, n1933, n1932}), .out(n583), .config_in(config_chain[4891:4890])); 
mux4 mux_141 (.in({n2545, n2544, n2535, n2534}), .out(n584), .config_in(config_chain[4893:4892])); 
mux4 mux_142 (.in({n1845, n1844, n1835, n1834}), .out(n585), .config_in(config_chain[4895:4894])); 
mux4 mux_143 (.in({n2445, n2444, n2435, n2434}), .out(n586), .config_in(config_chain[4897:4896])); 
mux4 mux_144 (.in({n1947, n1946, n1937, n1936}), .out(n587), .config_in(config_chain[4899:4898])); 
mux4 mux_145 (.in({n2547, n2546, n2537, n2536}), .out(n588), .config_in(config_chain[4901:4900])); 
mux4 mux_146 (.in({n1849, n1848, n1839, n1838}), .out(n589), .config_in(config_chain[4903:4902])); 
mux4 mux_147 (.in({n2449, n2448, n2439, n2438}), .out(n590), .config_in(config_chain[4905:4904])); 
mux4 mux_148 (.in({n2041, n2040, n2031, n2030}), .out(n609), .config_in(config_chain[4907:4906])); 
mux4 mux_149 (.in({n2561, n2560, n2551, n2550}), .out(n610), .config_in(config_chain[4909:4908])); 
mux4 mux_150 (.in({n1941, n1940, n1931, n1930}), .out(n611), .config_in(config_chain[4911:4910])); 
mux4 mux_151 (.in({n2463, n2462, n2453, n2452}), .out(n612), .config_in(config_chain[4913:4912])); 
mux4 mux_152 (.in({n2043, n2042, n2033, n2032}), .out(n613), .config_in(config_chain[4915:4914])); 
mux4 mux_153 (.in({n2565, n2564, n2555, n2554}), .out(n614), .config_in(config_chain[4917:4916])); 
mux4 mux_154 (.in({n1945, n1944, n1935, n1934}), .out(n615), .config_in(config_chain[4919:4918])); 
mux4 mux_155 (.in({n2465, n2464, n2455, n2454}), .out(n616), .config_in(config_chain[4921:4920])); 
mux4 mux_156 (.in({n2047, n2046, n2037, n2036}), .out(n617), .config_in(config_chain[4923:4922])); 
mux4 mux_157 (.in({n2567, n2566, n2557, n2556}), .out(n618), .config_in(config_chain[4925:4924])); 
mux4 mux_158 (.in({n1949, n1948, n1939, n1938}), .out(n619), .config_in(config_chain[4927:4926])); 
mux4 mux_159 (.in({n2469, n2468, n2459, n2458}), .out(n620), .config_in(config_chain[4929:4928])); 
mux4 mux_160 (.in({n2141, n2140, n2131, n2130}), .out(n639), .config_in(config_chain[4931:4930])); 
mux4 mux_161 (.in({n2581, n2580, n2571, n2570}), .out(n640), .config_in(config_chain[4933:4932])); 
mux4 mux_162 (.in({n2041, n2040, n2031, n2030}), .out(n641), .config_in(config_chain[4935:4934])); 
mux4 mux_163 (.in({n2483, n2482, n2473, n2472}), .out(n642), .config_in(config_chain[4937:4936])); 
mux4 mux_164 (.in({n2143, n2142, n2133, n2132}), .out(n643), .config_in(config_chain[4939:4938])); 
mux4 mux_165 (.in({n2585, n2584, n2575, n2574}), .out(n644), .config_in(config_chain[4941:4940])); 
mux4 mux_166 (.in({n2045, n2044, n2035, n2034}), .out(n645), .config_in(config_chain[4943:4942])); 
mux4 mux_167 (.in({n2485, n2484, n2475, n2474}), .out(n646), .config_in(config_chain[4945:4944])); 
mux4 mux_168 (.in({n2147, n2146, n2137, n2136}), .out(n647), .config_in(config_chain[4947:4946])); 
mux4 mux_169 (.in({n2587, n2586, n2577, n2576}), .out(n648), .config_in(config_chain[4949:4948])); 
mux4 mux_170 (.in({n2049, n2048, n2039, n2038}), .out(n649), .config_in(config_chain[4951:4950])); 
mux4 mux_171 (.in({n2489, n2488, n2479, n2478}), .out(n650), .config_in(config_chain[4953:4952])); 
mux4 mux_172 (.in({n2241, n2240, n2231, n2230}), .out(n669), .config_in(config_chain[4955:4954])); 
mux4 mux_173 (.in({n2601, n2600, n2591, n2590}), .out(n670), .config_in(config_chain[4957:4956])); 
mux4 mux_174 (.in({n2141, n2140, n2131, n2130}), .out(n671), .config_in(config_chain[4959:4958])); 
mux4 mux_175 (.in({n2503, n2502, n2493, n2492}), .out(n672), .config_in(config_chain[4961:4960])); 
mux4 mux_176 (.in({n2243, n2242, n2233, n2232}), .out(n673), .config_in(config_chain[4963:4962])); 
mux4 mux_177 (.in({n2605, n2604, n2595, n2594}), .out(n674), .config_in(config_chain[4965:4964])); 
mux4 mux_178 (.in({n2145, n2144, n2135, n2134}), .out(n675), .config_in(config_chain[4967:4966])); 
mux4 mux_179 (.in({n2505, n2504, n2495, n2494}), .out(n676), .config_in(config_chain[4969:4968])); 
mux4 mux_180 (.in({n2247, n2246, n2237, n2236}), .out(n677), .config_in(config_chain[4971:4970])); 
mux4 mux_181 (.in({n2607, n2606, n2597, n2596}), .out(n678), .config_in(config_chain[4973:4972])); 
mux4 mux_182 (.in({n2149, n2148, n2139, n2138}), .out(n679), .config_in(config_chain[4975:4974])); 
mux4 mux_183 (.in({n2509, n2508, n2499, n2498}), .out(n680), .config_in(config_chain[4977:4976])); 
mux4 mux_184 (.in({n2241, n2240, n2231, n2230}), .out(n708), .config_in(config_chain[4979:4978])); 
mux4 mux_185 (.in({n2241, n2240, n2231, n2230}), .out(n711), .config_in(config_chain[4981:4980])); 
mux4 mux_186 (.in({n2243, n2242, n2233, n2232}), .out(n714), .config_in(config_chain[4983:4982])); 
mux4 mux_187 (.in({n2245, n2244, n2235, n2234}), .out(n717), .config_in(config_chain[4985:4984])); 
mux4 mux_188 (.in({n2245, n2244, n2235, n2234}), .out(n720), .config_in(config_chain[4987:4986])); 
mux4 mux_189 (.in({n2247, n2246, n2237, n2236}), .out(n723), .config_in(config_chain[4989:4988])); 
mux4 mux_190 (.in({n2249, n2248, n2239, n2238}), .out(n726), .config_in(config_chain[4991:4990])); 
mux4 mux_191 (.in({n2249, n2248, n2239, n2238}), .out(n729), .config_in(config_chain[4993:4992])); 
mux4 mux_192 (.in({n1761, n1760, n1751, n1750}), .out(n756), .config_in(config_chain[4995:4994])); 
mux4 mux_193 (.in({n1761, n1760, n1751, n1750}), .out(n759), .config_in(config_chain[4997:4996])); 
mux4 mux_194 (.in({n1763, n1762, n1753, n1752}), .out(n762), .config_in(config_chain[4999:4998])); 
mux4 mux_195 (.in({n1763, n1762, n1753, n1752}), .out(n765), .config_in(config_chain[5001:5000])); 
mux4 mux_196 (.in({n1765, n1764, n1755, n1754}), .out(n768), .config_in(config_chain[5003:5002])); 
mux4 mux_197 (.in({n1767, n1766, n1757, n1756}), .out(n771), .config_in(config_chain[5005:5004])); 
mux4 mux_198 (.in({n1767, n1766, n1757, n1756}), .out(n774), .config_in(config_chain[5007:5006])); 
mux4 mux_199 (.in({n1769, n1768, n1759, n1758}), .out(n777), .config_in(config_chain[5009:5008])); 
mux4 mux_200 (.in({n1861, n1860, n1851, n1850}), .out(n795), .config_in(config_chain[5011:5010])); 
mux4 mux_201 (.in({n2621, n2620, n2611, n2610}), .out(n796), .config_in(config_chain[5013:5012])); 
mux4 mux_202 (.in({n1761, n1760, n1751, n1750}), .out(n797), .config_in(config_chain[5015:5014])); 
mux4 mux_203 (.in({n2523, n2522, n2513, n2512}), .out(n798), .config_in(config_chain[5017:5016])); 
mux4 mux_204 (.in({n1863, n1862, n1853, n1852}), .out(n799), .config_in(config_chain[5019:5018])); 
mux4 mux_205 (.in({n2625, n2624, n2615, n2614}), .out(n800), .config_in(config_chain[5021:5020])); 
mux4 mux_206 (.in({n1765, n1764, n1755, n1754}), .out(n801), .config_in(config_chain[5023:5022])); 
mux4 mux_207 (.in({n2525, n2524, n2515, n2514}), .out(n802), .config_in(config_chain[5025:5024])); 
mux4 mux_208 (.in({n1867, n1866, n1857, n1856}), .out(n803), .config_in(config_chain[5027:5026])); 
mux4 mux_209 (.in({n2627, n2626, n2617, n2616}), .out(n804), .config_in(config_chain[5029:5028])); 
mux4 mux_210 (.in({n1769, n1768, n1759, n1758}), .out(n805), .config_in(config_chain[5031:5030])); 
mux4 mux_211 (.in({n2529, n2528, n2519, n2518}), .out(n806), .config_in(config_chain[5033:5032])); 
mux4 mux_212 (.in({n1961, n1960, n1951, n1950}), .out(n825), .config_in(config_chain[5035:5034])); 
mux4 mux_213 (.in({n2641, n2640, n2631, n2630}), .out(n826), .config_in(config_chain[5037:5036])); 
mux4 mux_214 (.in({n1861, n1860, n1851, n1850}), .out(n827), .config_in(config_chain[5039:5038])); 
mux4 mux_215 (.in({n2543, n2542, n2533, n2532}), .out(n828), .config_in(config_chain[5041:5040])); 
mux4 mux_216 (.in({n1963, n1962, n1953, n1952}), .out(n829), .config_in(config_chain[5043:5042])); 
mux4 mux_217 (.in({n2645, n2644, n2635, n2634}), .out(n830), .config_in(config_chain[5045:5044])); 
mux4 mux_218 (.in({n1865, n1864, n1855, n1854}), .out(n831), .config_in(config_chain[5047:5046])); 
mux4 mux_219 (.in({n2545, n2544, n2535, n2534}), .out(n832), .config_in(config_chain[5049:5048])); 
mux4 mux_220 (.in({n1967, n1966, n1957, n1956}), .out(n833), .config_in(config_chain[5051:5050])); 
mux4 mux_221 (.in({n2647, n2646, n2637, n2636}), .out(n834), .config_in(config_chain[5053:5052])); 
mux4 mux_222 (.in({n1869, n1868, n1859, n1858}), .out(n835), .config_in(config_chain[5055:5054])); 
mux4 mux_223 (.in({n2549, n2548, n2539, n2538}), .out(n836), .config_in(config_chain[5057:5056])); 
mux4 mux_224 (.in({n2061, n2060, n2051, n2050}), .out(n855), .config_in(config_chain[5059:5058])); 
mux4 mux_225 (.in({n2661, n2660, n2651, n2650}), .out(n856), .config_in(config_chain[5061:5060])); 
mux4 mux_226 (.in({n1961, n1960, n1951, n1950}), .out(n857), .config_in(config_chain[5063:5062])); 
mux4 mux_227 (.in({n2563, n2562, n2553, n2552}), .out(n858), .config_in(config_chain[5065:5064])); 
mux4 mux_228 (.in({n2063, n2062, n2053, n2052}), .out(n859), .config_in(config_chain[5067:5066])); 
mux4 mux_229 (.in({n2665, n2664, n2655, n2654}), .out(n860), .config_in(config_chain[5069:5068])); 
mux4 mux_230 (.in({n1965, n1964, n1955, n1954}), .out(n861), .config_in(config_chain[5071:5070])); 
mux4 mux_231 (.in({n2565, n2564, n2555, n2554}), .out(n862), .config_in(config_chain[5073:5072])); 
mux4 mux_232 (.in({n2067, n2066, n2057, n2056}), .out(n863), .config_in(config_chain[5075:5074])); 
mux4 mux_233 (.in({n2667, n2666, n2657, n2656}), .out(n864), .config_in(config_chain[5077:5076])); 
mux4 mux_234 (.in({n1969, n1968, n1959, n1958}), .out(n865), .config_in(config_chain[5079:5078])); 
mux4 mux_235 (.in({n2569, n2568, n2559, n2558}), .out(n866), .config_in(config_chain[5081:5080])); 
mux4 mux_236 (.in({n2161, n2160, n2151, n2150}), .out(n885), .config_in(config_chain[5083:5082])); 
mux4 mux_237 (.in({n2681, n2680, n2671, n2670}), .out(n886), .config_in(config_chain[5085:5084])); 
mux4 mux_238 (.in({n2061, n2060, n2051, n2050}), .out(n887), .config_in(config_chain[5087:5086])); 
mux4 mux_239 (.in({n2583, n2582, n2573, n2572}), .out(n888), .config_in(config_chain[5089:5088])); 
mux4 mux_240 (.in({n2163, n2162, n2153, n2152}), .out(n889), .config_in(config_chain[5091:5090])); 
mux4 mux_241 (.in({n2685, n2684, n2675, n2674}), .out(n890), .config_in(config_chain[5093:5092])); 
mux4 mux_242 (.in({n2065, n2064, n2055, n2054}), .out(n891), .config_in(config_chain[5095:5094])); 
mux4 mux_243 (.in({n2585, n2584, n2575, n2574}), .out(n892), .config_in(config_chain[5097:5096])); 
mux4 mux_244 (.in({n2167, n2166, n2157, n2156}), .out(n893), .config_in(config_chain[5099:5098])); 
mux4 mux_245 (.in({n2687, n2686, n2677, n2676}), .out(n894), .config_in(config_chain[5101:5100])); 
mux4 mux_246 (.in({n2069, n2068, n2059, n2058}), .out(n895), .config_in(config_chain[5103:5102])); 
mux4 mux_247 (.in({n2589, n2588, n2579, n2578}), .out(n896), .config_in(config_chain[5105:5104])); 
mux4 mux_248 (.in({n2261, n2260, n2251, n2250}), .out(n915), .config_in(config_chain[5107:5106])); 
mux4 mux_249 (.in({n2701, n2700, n2691, n2690}), .out(n916), .config_in(config_chain[5109:5108])); 
mux4 mux_250 (.in({n2161, n2160, n2151, n2150}), .out(n917), .config_in(config_chain[5111:5110])); 
mux4 mux_251 (.in({n2603, n2602, n2593, n2592}), .out(n918), .config_in(config_chain[5113:5112])); 
mux4 mux_252 (.in({n2263, n2262, n2253, n2252}), .out(n919), .config_in(config_chain[5115:5114])); 
mux4 mux_253 (.in({n2705, n2704, n2695, n2694}), .out(n920), .config_in(config_chain[5117:5116])); 
mux4 mux_254 (.in({n2165, n2164, n2155, n2154}), .out(n921), .config_in(config_chain[5119:5118])); 
mux4 mux_255 (.in({n2605, n2604, n2595, n2594}), .out(n922), .config_in(config_chain[5121:5120])); 
mux4 mux_256 (.in({n2267, n2266, n2257, n2256}), .out(n923), .config_in(config_chain[5123:5122])); 
mux4 mux_257 (.in({n2707, n2706, n2697, n2696}), .out(n924), .config_in(config_chain[5125:5124])); 
mux4 mux_258 (.in({n2169, n2168, n2159, n2158}), .out(n925), .config_in(config_chain[5127:5126])); 
mux4 mux_259 (.in({n2609, n2608, n2599, n2598}), .out(n926), .config_in(config_chain[5129:5128])); 
mux4 mux_260 (.in({n2261, n2260, n2251, n2250}), .out(n954), .config_in(config_chain[5131:5130])); 
mux4 mux_261 (.in({n2261, n2260, n2251, n2250}), .out(n957), .config_in(config_chain[5133:5132])); 
mux4 mux_262 (.in({n2263, n2262, n2253, n2252}), .out(n960), .config_in(config_chain[5135:5134])); 
mux4 mux_263 (.in({n2265, n2264, n2255, n2254}), .out(n963), .config_in(config_chain[5137:5136])); 
mux4 mux_264 (.in({n2265, n2264, n2255, n2254}), .out(n966), .config_in(config_chain[5139:5138])); 
mux4 mux_265 (.in({n2267, n2266, n2257, n2256}), .out(n969), .config_in(config_chain[5141:5140])); 
mux4 mux_266 (.in({n2269, n2268, n2259, n2258}), .out(n972), .config_in(config_chain[5143:5142])); 
mux4 mux_267 (.in({n2269, n2268, n2259, n2258}), .out(n975), .config_in(config_chain[5145:5144])); 
mux4 mux_268 (.in({n1781, n1780, n1771, n1770}), .out(n1002), .config_in(config_chain[5147:5146])); 
mux4 mux_269 (.in({n1781, n1780, n1771, n1770}), .out(n1005), .config_in(config_chain[5149:5148])); 
mux4 mux_270 (.in({n1783, n1782, n1773, n1772}), .out(n1008), .config_in(config_chain[5151:5150])); 
mux4 mux_271 (.in({n1783, n1782, n1773, n1772}), .out(n1011), .config_in(config_chain[5153:5152])); 
mux4 mux_272 (.in({n1785, n1784, n1775, n1774}), .out(n1014), .config_in(config_chain[5155:5154])); 
mux4 mux_273 (.in({n1787, n1786, n1777, n1776}), .out(n1017), .config_in(config_chain[5157:5156])); 
mux4 mux_274 (.in({n1787, n1786, n1777, n1776}), .out(n1020), .config_in(config_chain[5159:5158])); 
mux4 mux_275 (.in({n1789, n1788, n1779, n1778}), .out(n1023), .config_in(config_chain[5161:5160])); 
mux4 mux_276 (.in({n1881, n1880, n1871, n1870}), .out(n1041), .config_in(config_chain[5163:5162])); 
mux4 mux_277 (.in({n2721, n2720, n2711, n2710}), .out(n1042), .config_in(config_chain[5165:5164])); 
mux4 mux_278 (.in({n1781, n1780, n1771, n1770}), .out(n1043), .config_in(config_chain[5167:5166])); 
mux4 mux_279 (.in({n2623, n2622, n2613, n2612}), .out(n1044), .config_in(config_chain[5169:5168])); 
mux4 mux_280 (.in({n1883, n1882, n1873, n1872}), .out(n1045), .config_in(config_chain[5171:5170])); 
mux4 mux_281 (.in({n2725, n2724, n2715, n2714}), .out(n1046), .config_in(config_chain[5173:5172])); 
mux4 mux_282 (.in({n1785, n1784, n1775, n1774}), .out(n1047), .config_in(config_chain[5175:5174])); 
mux4 mux_283 (.in({n2625, n2624, n2615, n2614}), .out(n1048), .config_in(config_chain[5177:5176])); 
mux4 mux_284 (.in({n1887, n1886, n1877, n1876}), .out(n1049), .config_in(config_chain[5179:5178])); 
mux4 mux_285 (.in({n2727, n2726, n2717, n2716}), .out(n1050), .config_in(config_chain[5181:5180])); 
mux4 mux_286 (.in({n1789, n1788, n1779, n1778}), .out(n1051), .config_in(config_chain[5183:5182])); 
mux4 mux_287 (.in({n2629, n2628, n2619, n2618}), .out(n1052), .config_in(config_chain[5185:5184])); 
mux4 mux_288 (.in({n1981, n1980, n1971, n1970}), .out(n1071), .config_in(config_chain[5187:5186])); 
mux4 mux_289 (.in({n2741, n2740, n2731, n2730}), .out(n1072), .config_in(config_chain[5189:5188])); 
mux4 mux_290 (.in({n1881, n1880, n1871, n1870}), .out(n1073), .config_in(config_chain[5191:5190])); 
mux4 mux_291 (.in({n2643, n2642, n2633, n2632}), .out(n1074), .config_in(config_chain[5193:5192])); 
mux4 mux_292 (.in({n1983, n1982, n1973, n1972}), .out(n1075), .config_in(config_chain[5195:5194])); 
mux4 mux_293 (.in({n2745, n2744, n2735, n2734}), .out(n1076), .config_in(config_chain[5197:5196])); 
mux4 mux_294 (.in({n1885, n1884, n1875, n1874}), .out(n1077), .config_in(config_chain[5199:5198])); 
mux4 mux_295 (.in({n2645, n2644, n2635, n2634}), .out(n1078), .config_in(config_chain[5201:5200])); 
mux4 mux_296 (.in({n1987, n1986, n1977, n1976}), .out(n1079), .config_in(config_chain[5203:5202])); 
mux4 mux_297 (.in({n2747, n2746, n2737, n2736}), .out(n1080), .config_in(config_chain[5205:5204])); 
mux4 mux_298 (.in({n1889, n1888, n1879, n1878}), .out(n1081), .config_in(config_chain[5207:5206])); 
mux4 mux_299 (.in({n2649, n2648, n2639, n2638}), .out(n1082), .config_in(config_chain[5209:5208])); 
mux4 mux_300 (.in({n2081, n2080, n2071, n2070}), .out(n1101), .config_in(config_chain[5211:5210])); 
mux4 mux_301 (.in({n2761, n2760, n2751, n2750}), .out(n1102), .config_in(config_chain[5213:5212])); 
mux4 mux_302 (.in({n1981, n1980, n1971, n1970}), .out(n1103), .config_in(config_chain[5215:5214])); 
mux4 mux_303 (.in({n2663, n2662, n2653, n2652}), .out(n1104), .config_in(config_chain[5217:5216])); 
mux4 mux_304 (.in({n2083, n2082, n2073, n2072}), .out(n1105), .config_in(config_chain[5219:5218])); 
mux4 mux_305 (.in({n2765, n2764, n2755, n2754}), .out(n1106), .config_in(config_chain[5221:5220])); 
mux4 mux_306 (.in({n1985, n1984, n1975, n1974}), .out(n1107), .config_in(config_chain[5223:5222])); 
mux4 mux_307 (.in({n2665, n2664, n2655, n2654}), .out(n1108), .config_in(config_chain[5225:5224])); 
mux4 mux_308 (.in({n2087, n2086, n2077, n2076}), .out(n1109), .config_in(config_chain[5227:5226])); 
mux4 mux_309 (.in({n2767, n2766, n2757, n2756}), .out(n1110), .config_in(config_chain[5229:5228])); 
mux4 mux_310 (.in({n1989, n1988, n1979, n1978}), .out(n1111), .config_in(config_chain[5231:5230])); 
mux4 mux_311 (.in({n2669, n2668, n2659, n2658}), .out(n1112), .config_in(config_chain[5233:5232])); 
mux4 mux_312 (.in({n2181, n2180, n2171, n2170}), .out(n1131), .config_in(config_chain[5235:5234])); 
mux4 mux_313 (.in({n2781, n2780, n2771, n2770}), .out(n1132), .config_in(config_chain[5237:5236])); 
mux4 mux_314 (.in({n2081, n2080, n2071, n2070}), .out(n1133), .config_in(config_chain[5239:5238])); 
mux4 mux_315 (.in({n2683, n2682, n2673, n2672}), .out(n1134), .config_in(config_chain[5241:5240])); 
mux4 mux_316 (.in({n2183, n2182, n2173, n2172}), .out(n1135), .config_in(config_chain[5243:5242])); 
mux4 mux_317 (.in({n2785, n2784, n2775, n2774}), .out(n1136), .config_in(config_chain[5245:5244])); 
mux4 mux_318 (.in({n2085, n2084, n2075, n2074}), .out(n1137), .config_in(config_chain[5247:5246])); 
mux4 mux_319 (.in({n2685, n2684, n2675, n2674}), .out(n1138), .config_in(config_chain[5249:5248])); 
mux4 mux_320 (.in({n2187, n2186, n2177, n2176}), .out(n1139), .config_in(config_chain[5251:5250])); 
mux4 mux_321 (.in({n2787, n2786, n2777, n2776}), .out(n1140), .config_in(config_chain[5253:5252])); 
mux4 mux_322 (.in({n2089, n2088, n2079, n2078}), .out(n1141), .config_in(config_chain[5255:5254])); 
mux4 mux_323 (.in({n2689, n2688, n2679, n2678}), .out(n1142), .config_in(config_chain[5257:5256])); 
mux4 mux_324 (.in({n2281, n2280, n2271, n2270}), .out(n1161), .config_in(config_chain[5259:5258])); 
mux4 mux_325 (.in({n2801, n2800, n2791, n2790}), .out(n1162), .config_in(config_chain[5261:5260])); 
mux4 mux_326 (.in({n2181, n2180, n2171, n2170}), .out(n1163), .config_in(config_chain[5263:5262])); 
mux4 mux_327 (.in({n2703, n2702, n2693, n2692}), .out(n1164), .config_in(config_chain[5265:5264])); 
mux4 mux_328 (.in({n2283, n2282, n2273, n2272}), .out(n1165), .config_in(config_chain[5267:5266])); 
mux4 mux_329 (.in({n2805, n2804, n2795, n2794}), .out(n1166), .config_in(config_chain[5269:5268])); 
mux4 mux_330 (.in({n2185, n2184, n2175, n2174}), .out(n1167), .config_in(config_chain[5271:5270])); 
mux4 mux_331 (.in({n2705, n2704, n2695, n2694}), .out(n1168), .config_in(config_chain[5273:5272])); 
mux4 mux_332 (.in({n2287, n2286, n2277, n2276}), .out(n1169), .config_in(config_chain[5275:5274])); 
mux4 mux_333 (.in({n2807, n2806, n2797, n2796}), .out(n1170), .config_in(config_chain[5277:5276])); 
mux4 mux_334 (.in({n2189, n2188, n2179, n2178}), .out(n1171), .config_in(config_chain[5279:5278])); 
mux4 mux_335 (.in({n2709, n2708, n2699, n2698}), .out(n1172), .config_in(config_chain[5281:5280])); 
mux4 mux_336 (.in({n2281, n2280, n2271, n2270}), .out(n1200), .config_in(config_chain[5283:5282])); 
mux4 mux_337 (.in({n2281, n2280, n2271, n2270}), .out(n1203), .config_in(config_chain[5285:5284])); 
mux4 mux_338 (.in({n2283, n2282, n2273, n2272}), .out(n1206), .config_in(config_chain[5287:5286])); 
mux4 mux_339 (.in({n2285, n2284, n2275, n2274}), .out(n1209), .config_in(config_chain[5289:5288])); 
mux4 mux_340 (.in({n2285, n2284, n2275, n2274}), .out(n1212), .config_in(config_chain[5291:5290])); 
mux4 mux_341 (.in({n2287, n2286, n2277, n2276}), .out(n1215), .config_in(config_chain[5293:5292])); 
mux4 mux_342 (.in({n2289, n2288, n2279, n2278}), .out(n1218), .config_in(config_chain[5295:5294])); 
mux4 mux_343 (.in({n2289, n2288, n2279, n2278}), .out(n1221), .config_in(config_chain[5297:5296])); 
mux4 mux_344 (.in({n1801, n1800, n1791, n1790}), .out(n1248), .config_in(config_chain[5299:5298])); 
mux4 mux_345 (.in({n1801, n1800, n1791, n1790}), .out(n1251), .config_in(config_chain[5301:5300])); 
mux4 mux_346 (.in({n1803, n1802, n1793, n1792}), .out(n1254), .config_in(config_chain[5303:5302])); 
mux4 mux_347 (.in({n1803, n1802, n1793, n1792}), .out(n1257), .config_in(config_chain[5305:5304])); 
mux4 mux_348 (.in({n1805, n1804, n1795, n1794}), .out(n1260), .config_in(config_chain[5307:5306])); 
mux4 mux_349 (.in({n1807, n1806, n1797, n1796}), .out(n1263), .config_in(config_chain[5309:5308])); 
mux4 mux_350 (.in({n1807, n1806, n1797, n1796}), .out(n1266), .config_in(config_chain[5311:5310])); 
mux4 mux_351 (.in({n1809, n1808, n1799, n1798}), .out(n1269), .config_in(config_chain[5313:5312])); 
mux4 mux_352 (.in({n1901, n1900, n1891, n1890}), .out(n1287), .config_in(config_chain[5315:5314])); 
mux4 mux_353 (.in({n2821, n2820, n2811, n2810}), .out(n1288), .config_in(config_chain[5317:5316])); 
mux4 mux_354 (.in({n1801, n1800, n1791, n1790}), .out(n1289), .config_in(config_chain[5319:5318])); 
mux4 mux_355 (.in({n2723, n2722, n2713, n2712}), .out(n1290), .config_in(config_chain[5321:5320])); 
mux4 mux_356 (.in({n1903, n1902, n1893, n1892}), .out(n1291), .config_in(config_chain[5323:5322])); 
mux4 mux_357 (.in({n2825, n2824, n2815, n2814}), .out(n1292), .config_in(config_chain[5325:5324])); 
mux4 mux_358 (.in({n1805, n1804, n1795, n1794}), .out(n1293), .config_in(config_chain[5327:5326])); 
mux4 mux_359 (.in({n2725, n2724, n2715, n2714}), .out(n1294), .config_in(config_chain[5329:5328])); 
mux4 mux_360 (.in({n1907, n1906, n1897, n1896}), .out(n1295), .config_in(config_chain[5331:5330])); 
mux4 mux_361 (.in({n2827, n2826, n2817, n2816}), .out(n1296), .config_in(config_chain[5333:5332])); 
mux4 mux_362 (.in({n1809, n1808, n1799, n1798}), .out(n1297), .config_in(config_chain[5335:5334])); 
mux4 mux_363 (.in({n2729, n2728, n2719, n2718}), .out(n1298), .config_in(config_chain[5337:5336])); 
mux4 mux_364 (.in({n2001, n2000, n1991, n1990}), .out(n1317), .config_in(config_chain[5339:5338])); 
mux4 mux_365 (.in({n2841, n2840, n2831, n2830}), .out(n1318), .config_in(config_chain[5341:5340])); 
mux4 mux_366 (.in({n1901, n1900, n1891, n1890}), .out(n1319), .config_in(config_chain[5343:5342])); 
mux4 mux_367 (.in({n2743, n2742, n2733, n2732}), .out(n1320), .config_in(config_chain[5345:5344])); 
mux4 mux_368 (.in({n2003, n2002, n1993, n1992}), .out(n1321), .config_in(config_chain[5347:5346])); 
mux4 mux_369 (.in({n2845, n2844, n2835, n2834}), .out(n1322), .config_in(config_chain[5349:5348])); 
mux4 mux_370 (.in({n1905, n1904, n1895, n1894}), .out(n1323), .config_in(config_chain[5351:5350])); 
mux4 mux_371 (.in({n2745, n2744, n2735, n2734}), .out(n1324), .config_in(config_chain[5353:5352])); 
mux4 mux_372 (.in({n2007, n2006, n1997, n1996}), .out(n1325), .config_in(config_chain[5355:5354])); 
mux4 mux_373 (.in({n2847, n2846, n2837, n2836}), .out(n1326), .config_in(config_chain[5357:5356])); 
mux4 mux_374 (.in({n1909, n1908, n1899, n1898}), .out(n1327), .config_in(config_chain[5359:5358])); 
mux4 mux_375 (.in({n2749, n2748, n2739, n2738}), .out(n1328), .config_in(config_chain[5361:5360])); 
mux4 mux_376 (.in({n2101, n2100, n2091, n2090}), .out(n1347), .config_in(config_chain[5363:5362])); 
mux4 mux_377 (.in({n2861, n2860, n2851, n2850}), .out(n1348), .config_in(config_chain[5365:5364])); 
mux4 mux_378 (.in({n2001, n2000, n1991, n1990}), .out(n1349), .config_in(config_chain[5367:5366])); 
mux4 mux_379 (.in({n2763, n2762, n2753, n2752}), .out(n1350), .config_in(config_chain[5369:5368])); 
mux4 mux_380 (.in({n2103, n2102, n2093, n2092}), .out(n1351), .config_in(config_chain[5371:5370])); 
mux4 mux_381 (.in({n2865, n2864, n2855, n2854}), .out(n1352), .config_in(config_chain[5373:5372])); 
mux4 mux_382 (.in({n2005, n2004, n1995, n1994}), .out(n1353), .config_in(config_chain[5375:5374])); 
mux4 mux_383 (.in({n2765, n2764, n2755, n2754}), .out(n1354), .config_in(config_chain[5377:5376])); 
mux4 mux_384 (.in({n2107, n2106, n2097, n2096}), .out(n1355), .config_in(config_chain[5379:5378])); 
mux4 mux_385 (.in({n2867, n2866, n2857, n2856}), .out(n1356), .config_in(config_chain[5381:5380])); 
mux4 mux_386 (.in({n2009, n2008, n1999, n1998}), .out(n1357), .config_in(config_chain[5383:5382])); 
mux4 mux_387 (.in({n2769, n2768, n2759, n2758}), .out(n1358), .config_in(config_chain[5385:5384])); 
mux4 mux_388 (.in({n2201, n2200, n2191, n2190}), .out(n1377), .config_in(config_chain[5387:5386])); 
mux4 mux_389 (.in({n2881, n2880, n2871, n2870}), .out(n1378), .config_in(config_chain[5389:5388])); 
mux4 mux_390 (.in({n2101, n2100, n2091, n2090}), .out(n1379), .config_in(config_chain[5391:5390])); 
mux4 mux_391 (.in({n2783, n2782, n2773, n2772}), .out(n1380), .config_in(config_chain[5393:5392])); 
mux4 mux_392 (.in({n2203, n2202, n2193, n2192}), .out(n1381), .config_in(config_chain[5395:5394])); 
mux4 mux_393 (.in({n2885, n2884, n2875, n2874}), .out(n1382), .config_in(config_chain[5397:5396])); 
mux4 mux_394 (.in({n2105, n2104, n2095, n2094}), .out(n1383), .config_in(config_chain[5399:5398])); 
mux4 mux_395 (.in({n2785, n2784, n2775, n2774}), .out(n1384), .config_in(config_chain[5401:5400])); 
mux4 mux_396 (.in({n2207, n2206, n2197, n2196}), .out(n1385), .config_in(config_chain[5403:5402])); 
mux4 mux_397 (.in({n2887, n2886, n2877, n2876}), .out(n1386), .config_in(config_chain[5405:5404])); 
mux4 mux_398 (.in({n2109, n2108, n2099, n2098}), .out(n1387), .config_in(config_chain[5407:5406])); 
mux4 mux_399 (.in({n2789, n2788, n2779, n2778}), .out(n1388), .config_in(config_chain[5409:5408])); 
mux4 mux_400 (.in({n2301, n2300, n2291, n2290}), .out(n1407), .config_in(config_chain[5411:5410])); 
mux4 mux_401 (.in({n2901, n2900, n2891, n2890}), .out(n1408), .config_in(config_chain[5413:5412])); 
mux4 mux_402 (.in({n2201, n2200, n2191, n2190}), .out(n1409), .config_in(config_chain[5415:5414])); 
mux4 mux_403 (.in({n2803, n2802, n2793, n2792}), .out(n1410), .config_in(config_chain[5417:5416])); 
mux4 mux_404 (.in({n2303, n2302, n2293, n2292}), .out(n1411), .config_in(config_chain[5419:5418])); 
mux4 mux_405 (.in({n2905, n2904, n2895, n2894}), .out(n1412), .config_in(config_chain[5421:5420])); 
mux4 mux_406 (.in({n2205, n2204, n2195, n2194}), .out(n1413), .config_in(config_chain[5423:5422])); 
mux4 mux_407 (.in({n2805, n2804, n2795, n2794}), .out(n1414), .config_in(config_chain[5425:5424])); 
mux4 mux_408 (.in({n2307, n2306, n2297, n2296}), .out(n1415), .config_in(config_chain[5427:5426])); 
mux4 mux_409 (.in({n2907, n2906, n2897, n2896}), .out(n1416), .config_in(config_chain[5429:5428])); 
mux4 mux_410 (.in({n2209, n2208, n2199, n2198}), .out(n1417), .config_in(config_chain[5431:5430])); 
mux4 mux_411 (.in({n2809, n2808, n2799, n2798}), .out(n1418), .config_in(config_chain[5433:5432])); 
mux4 mux_412 (.in({n2301, n2300, n2291, n2290}), .out(n1446), .config_in(config_chain[5435:5434])); 
mux4 mux_413 (.in({n2301, n2300, n2291, n2290}), .out(n1449), .config_in(config_chain[5437:5436])); 
mux4 mux_414 (.in({n2303, n2302, n2293, n2292}), .out(n1452), .config_in(config_chain[5439:5438])); 
mux4 mux_415 (.in({n2305, n2304, n2295, n2294}), .out(n1455), .config_in(config_chain[5441:5440])); 
mux4 mux_416 (.in({n2305, n2304, n2295, n2294}), .out(n1458), .config_in(config_chain[5443:5442])); 
mux4 mux_417 (.in({n2307, n2306, n2297, n2296}), .out(n1461), .config_in(config_chain[5445:5444])); 
mux4 mux_418 (.in({n2309, n2308, n2299, n2298}), .out(n1464), .config_in(config_chain[5447:5446])); 
mux4 mux_419 (.in({n2309, n2308, n2299, n2298}), .out(n1467), .config_in(config_chain[5449:5448])); 
mux4 mux_420 (.in({n2821, n2820, n2811, n2810}), .out(n1494), .config_in(config_chain[5451:5450])); 
mux4 mux_421 (.in({n2823, n2822, n2813, n2812}), .out(n1497), .config_in(config_chain[5453:5452])); 
mux4 mux_422 (.in({n2823, n2822, n2813, n2812}), .out(n1500), .config_in(config_chain[5455:5454])); 
mux4 mux_423 (.in({n2825, n2824, n2815, n2814}), .out(n1503), .config_in(config_chain[5457:5456])); 
mux4 mux_424 (.in({n2825, n2824, n2815, n2814}), .out(n1506), .config_in(config_chain[5459:5458])); 
mux4 mux_425 (.in({n2827, n2826, n2817, n2816}), .out(n1509), .config_in(config_chain[5461:5460])); 
mux4 mux_426 (.in({n2829, n2828, n2819, n2818}), .out(n1512), .config_in(config_chain[5463:5462])); 
mux4 mux_427 (.in({n2829, n2828, n2819, n2818}), .out(n1515), .config_in(config_chain[5465:5464])); 
mux4 mux_428 (.in({n2841, n2840, n2831, n2830}), .out(n1542), .config_in(config_chain[5467:5466])); 
mux4 mux_429 (.in({n2843, n2842, n2833, n2832}), .out(n1545), .config_in(config_chain[5469:5468])); 
mux4 mux_430 (.in({n2843, n2842, n2833, n2832}), .out(n1548), .config_in(config_chain[5471:5470])); 
mux4 mux_431 (.in({n2845, n2844, n2835, n2834}), .out(n1551), .config_in(config_chain[5473:5472])); 
mux4 mux_432 (.in({n2845, n2844, n2835, n2834}), .out(n1554), .config_in(config_chain[5475:5474])); 
mux4 mux_433 (.in({n2847, n2846, n2837, n2836}), .out(n1557), .config_in(config_chain[5477:5476])); 
mux4 mux_434 (.in({n2849, n2848, n2839, n2838}), .out(n1560), .config_in(config_chain[5479:5478])); 
mux4 mux_435 (.in({n2849, n2848, n2839, n2838}), .out(n1563), .config_in(config_chain[5481:5480])); 
mux4 mux_436 (.in({n2861, n2860, n2851, n2850}), .out(n1590), .config_in(config_chain[5483:5482])); 
mux4 mux_437 (.in({n2863, n2862, n2853, n2852}), .out(n1593), .config_in(config_chain[5485:5484])); 
mux4 mux_438 (.in({n2863, n2862, n2853, n2852}), .out(n1596), .config_in(config_chain[5487:5486])); 
mux4 mux_439 (.in({n2865, n2864, n2855, n2854}), .out(n1599), .config_in(config_chain[5489:5488])); 
mux4 mux_440 (.in({n2865, n2864, n2855, n2854}), .out(n1602), .config_in(config_chain[5491:5490])); 
mux4 mux_441 (.in({n2867, n2866, n2857, n2856}), .out(n1605), .config_in(config_chain[5493:5492])); 
mux4 mux_442 (.in({n2869, n2868, n2859, n2858}), .out(n1608), .config_in(config_chain[5495:5494])); 
mux4 mux_443 (.in({n2869, n2868, n2859, n2858}), .out(n1611), .config_in(config_chain[5497:5496])); 
mux4 mux_444 (.in({n2881, n2880, n2871, n2870}), .out(n1638), .config_in(config_chain[5499:5498])); 
mux4 mux_445 (.in({n2883, n2882, n2873, n2872}), .out(n1641), .config_in(config_chain[5501:5500])); 
mux4 mux_446 (.in({n2883, n2882, n2873, n2872}), .out(n1644), .config_in(config_chain[5503:5502])); 
mux4 mux_447 (.in({n2885, n2884, n2875, n2874}), .out(n1647), .config_in(config_chain[5505:5504])); 
mux4 mux_448 (.in({n2885, n2884, n2875, n2874}), .out(n1650), .config_in(config_chain[5507:5506])); 
mux4 mux_449 (.in({n2887, n2886, n2877, n2876}), .out(n1653), .config_in(config_chain[5509:5508])); 
mux4 mux_450 (.in({n2889, n2888, n2879, n2878}), .out(n1656), .config_in(config_chain[5511:5510])); 
mux4 mux_451 (.in({n2889, n2888, n2879, n2878}), .out(n1659), .config_in(config_chain[5513:5512])); 
mux4 mux_452 (.in({n2901, n2900, n2891, n2890}), .out(n1686), .config_in(config_chain[5515:5514])); 
mux4 mux_453 (.in({n2903, n2902, n2893, n2892}), .out(n1689), .config_in(config_chain[5517:5516])); 
mux4 mux_454 (.in({n2903, n2902, n2893, n2892}), .out(n1692), .config_in(config_chain[5519:5518])); 
mux4 mux_455 (.in({n2905, n2904, n2895, n2894}), .out(n1695), .config_in(config_chain[5521:5520])); 
mux4 mux_456 (.in({n2905, n2904, n2895, n2894}), .out(n1698), .config_in(config_chain[5523:5522])); 
mux4 mux_457 (.in({n2907, n2906, n2897, n2896}), .out(n1701), .config_in(config_chain[5525:5524])); 
mux4 mux_458 (.in({n2909, n2908, n2899, n2898}), .out(n1704), .config_in(config_chain[5527:5526])); 
mux4 mux_459 (.in({n2909, n2908, n2899, n2898}), .out(n1707), .config_in(config_chain[5529:5528])); 
mux3 mux_460 (.in({n2329, n280, n265}), .out(n1710), .config_in(config_chain[5531:5530])); 
mux4 mux_461 (.in({n2411, n1731, n280, n265}), .out(n1711), .config_in(config_chain[5533:5532])); 
mux3 mux_462 (.in({n2311, n280, n265}), .out(n1712), .config_in(config_chain[5535:5534])); 
mux4 mux_463 (.in({n2413, n1733, n280, n265}), .out(n1713), .config_in(config_chain[5537:5536])); 
mux3 mux_464 (.in({n2313, n283, n268}), .out(n1714), .config_in(config_chain[5539:5538])); 
mux4 mux_465 (.in({n2415, n1735, n283, n268}), .out(n1715), .config_in(config_chain[5541:5540])); 
mux3 mux_466 (.in({n2315, n283, n268}), .out(n1716), .config_in(config_chain[5543:5542])); 
mux4 mux_467 (.in({n2417, n1737, n283, n268}), .out(n1717), .config_in(config_chain[5545:5544])); 
mux3 mux_468 (.in({n2317, n286, n271}), .out(n1718), .config_in(config_chain[5547:5546])); 
mux4 mux_469 (.in({n2419, n1739, n286, n271}), .out(n1719), .config_in(config_chain[5549:5548])); 
mux3 mux_470 (.in({n2319, n286, n271}), .out(n1720), .config_in(config_chain[5551:5550])); 
mux4 mux_471 (.in({n2421, n1741, n286, n271}), .out(n1721), .config_in(config_chain[5553:5552])); 
mux2 mux_472 (.in({n2321, n274}), .out(n1722), .config_in(config_chain[5554:5554])); 
mux3 mux_473 (.in({n2423, n1743, n274}), .out(n1723), .config_in(config_chain[5556:5555])); 
mux2 mux_474 (.in({n2323, n274}), .out(n1724), .config_in(config_chain[5557:5557])); 
mux3 mux_475 (.in({n2425, n1745, n274}), .out(n1725), .config_in(config_chain[5559:5558])); 
mux2 mux_476 (.in({n2325, n277}), .out(n1726), .config_in(config_chain[5560:5560])); 
mux3 mux_477 (.in({n2427, n1747, n277}), .out(n1727), .config_in(config_chain[5562:5561])); 
mux2 mux_478 (.in({n2327, n277}), .out(n1728), .config_in(config_chain[5563:5563])); 
mux3 mux_479 (.in({n2429, n1749, n277}), .out(n1729), .config_in(config_chain[5565:5564])); 
mux4 mux_480 (.in({n2411, n1710, n526, n511}), .out(n1730), .config_in(config_chain[5567:5566])); 
mux4 mux_481 (.in({n2511, n1751, n526, n511}), .out(n1731), .config_in(config_chain[5569:5568])); 
mux4 mux_482 (.in({n2413, n1712, n526, n511}), .out(n1732), .config_in(config_chain[5571:5570])); 
mux4 mux_483 (.in({n2513, n1753, n526, n511}), .out(n1733), .config_in(config_chain[5573:5572])); 
mux4 mux_484 (.in({n2415, n1714, n529, n514}), .out(n1734), .config_in(config_chain[5575:5574])); 
mux4 mux_485 (.in({n2515, n1755, n529, n514}), .out(n1735), .config_in(config_chain[5577:5576])); 
mux4 mux_486 (.in({n2417, n1716, n529, n514}), .out(n1736), .config_in(config_chain[5579:5578])); 
mux4 mux_487 (.in({n2517, n1757, n529, n514}), .out(n1737), .config_in(config_chain[5581:5580])); 
mux4 mux_488 (.in({n2419, n1718, n532, n517}), .out(n1738), .config_in(config_chain[5583:5582])); 
mux4 mux_489 (.in({n2519, n1759, n532, n517}), .out(n1739), .config_in(config_chain[5585:5584])); 
mux4 mux_490 (.in({n2421, n1720, n532, n517}), .out(n1740), .config_in(config_chain[5587:5586])); 
mux4 mux_491 (.in({n2521, n1761, n532, n517}), .out(n1741), .config_in(config_chain[5589:5588])); 
mux3 mux_492 (.in({n2423, n1722, n520}), .out(n1742), .config_in(config_chain[5591:5590])); 
mux3 mux_493 (.in({n2523, n1763, n520}), .out(n1743), .config_in(config_chain[5593:5592])); 
mux3 mux_494 (.in({n2425, n1724, n520}), .out(n1744), .config_in(config_chain[5595:5594])); 
mux3 mux_495 (.in({n2525, n1765, n520}), .out(n1745), .config_in(config_chain[5597:5596])); 
mux3 mux_496 (.in({n2427, n1726, n523}), .out(n1746), .config_in(config_chain[5599:5598])); 
mux3 mux_497 (.in({n2527, n1767, n523}), .out(n1747), .config_in(config_chain[5601:5600])); 
mux3 mux_498 (.in({n2429, n1728, n523}), .out(n1748), .config_in(config_chain[5603:5602])); 
mux3 mux_499 (.in({n2529, n1769, n523}), .out(n1749), .config_in(config_chain[5605:5604])); 
mux4 mux_500 (.in({n2511, n1730, n772, n757}), .out(n1750), .config_in(config_chain[5607:5606])); 
mux4 mux_501 (.in({n2611, n1771, n772, n757}), .out(n1751), .config_in(config_chain[5609:5608])); 
mux4 mux_502 (.in({n2513, n1732, n772, n757}), .out(n1752), .config_in(config_chain[5611:5610])); 
mux4 mux_503 (.in({n2613, n1773, n772, n757}), .out(n1753), .config_in(config_chain[5613:5612])); 
mux4 mux_504 (.in({n2515, n1734, n775, n760}), .out(n1754), .config_in(config_chain[5615:5614])); 
mux4 mux_505 (.in({n2615, n1775, n775, n760}), .out(n1755), .config_in(config_chain[5617:5616])); 
mux4 mux_506 (.in({n2517, n1736, n775, n760}), .out(n1756), .config_in(config_chain[5619:5618])); 
mux4 mux_507 (.in({n2617, n1777, n775, n760}), .out(n1757), .config_in(config_chain[5621:5620])); 
mux4 mux_508 (.in({n2519, n1738, n778, n763}), .out(n1758), .config_in(config_chain[5623:5622])); 
mux4 mux_509 (.in({n2619, n1779, n778, n763}), .out(n1759), .config_in(config_chain[5625:5624])); 
mux4 mux_510 (.in({n2521, n1740, n778, n763}), .out(n1760), .config_in(config_chain[5627:5626])); 
mux4 mux_511 (.in({n2621, n1781, n778, n763}), .out(n1761), .config_in(config_chain[5629:5628])); 
mux3 mux_512 (.in({n2523, n1742, n766}), .out(n1762), .config_in(config_chain[5631:5630])); 
mux3 mux_513 (.in({n2623, n1783, n766}), .out(n1763), .config_in(config_chain[5633:5632])); 
mux3 mux_514 (.in({n2525, n1744, n766}), .out(n1764), .config_in(config_chain[5635:5634])); 
mux3 mux_515 (.in({n2625, n1785, n766}), .out(n1765), .config_in(config_chain[5637:5636])); 
mux3 mux_516 (.in({n2527, n1746, n769}), .out(n1766), .config_in(config_chain[5639:5638])); 
mux3 mux_517 (.in({n2627, n1787, n769}), .out(n1767), .config_in(config_chain[5641:5640])); 
mux3 mux_518 (.in({n2529, n1748, n769}), .out(n1768), .config_in(config_chain[5643:5642])); 
mux3 mux_519 (.in({n2629, n1789, n769}), .out(n1769), .config_in(config_chain[5645:5644])); 
mux4 mux_520 (.in({n2611, n1750, n1018, n1003}), .out(n1770), .config_in(config_chain[5647:5646])); 
mux4 mux_521 (.in({n2711, n1791, n1018, n1003}), .out(n1771), .config_in(config_chain[5649:5648])); 
mux4 mux_522 (.in({n2613, n1752, n1018, n1003}), .out(n1772), .config_in(config_chain[5651:5650])); 
mux4 mux_523 (.in({n2713, n1793, n1018, n1003}), .out(n1773), .config_in(config_chain[5653:5652])); 
mux4 mux_524 (.in({n2615, n1754, n1021, n1006}), .out(n1774), .config_in(config_chain[5655:5654])); 
mux4 mux_525 (.in({n2715, n1795, n1021, n1006}), .out(n1775), .config_in(config_chain[5657:5656])); 
mux4 mux_526 (.in({n2617, n1756, n1021, n1006}), .out(n1776), .config_in(config_chain[5659:5658])); 
mux4 mux_527 (.in({n2717, n1797, n1021, n1006}), .out(n1777), .config_in(config_chain[5661:5660])); 
mux4 mux_528 (.in({n2619, n1758, n1024, n1009}), .out(n1778), .config_in(config_chain[5663:5662])); 
mux4 mux_529 (.in({n2719, n1799, n1024, n1009}), .out(n1779), .config_in(config_chain[5665:5664])); 
mux4 mux_530 (.in({n2621, n1760, n1024, n1009}), .out(n1780), .config_in(config_chain[5667:5666])); 
mux4 mux_531 (.in({n2721, n1801, n1024, n1009}), .out(n1781), .config_in(config_chain[5669:5668])); 
mux3 mux_532 (.in({n2623, n1762, n1012}), .out(n1782), .config_in(config_chain[5671:5670])); 
mux3 mux_533 (.in({n2723, n1803, n1012}), .out(n1783), .config_in(config_chain[5673:5672])); 
mux3 mux_534 (.in({n2625, n1764, n1012}), .out(n1784), .config_in(config_chain[5675:5674])); 
mux3 mux_535 (.in({n2725, n1805, n1012}), .out(n1785), .config_in(config_chain[5677:5676])); 
mux3 mux_536 (.in({n2627, n1766, n1015}), .out(n1786), .config_in(config_chain[5679:5678])); 
mux3 mux_537 (.in({n2727, n1807, n1015}), .out(n1787), .config_in(config_chain[5681:5680])); 
mux3 mux_538 (.in({n2629, n1768, n1015}), .out(n1788), .config_in(config_chain[5683:5682])); 
mux3 mux_539 (.in({n2729, n1809, n1015}), .out(n1789), .config_in(config_chain[5685:5684])); 
mux4 mux_540 (.in({n2711, n1770, n1264, n1249}), .out(n1790), .config_in(config_chain[5687:5686])); 
mux3 mux_541 (.in({n2811, n1264, n1249}), .out(n1791), .config_in(config_chain[5689:5688])); 
mux4 mux_542 (.in({n2713, n1772, n1264, n1249}), .out(n1792), .config_in(config_chain[5691:5690])); 
mux3 mux_543 (.in({n2829, n1264, n1249}), .out(n1793), .config_in(config_chain[5693:5692])); 
mux4 mux_544 (.in({n2715, n1774, n1267, n1252}), .out(n1794), .config_in(config_chain[5695:5694])); 
mux3 mux_545 (.in({n2827, n1267, n1252}), .out(n1795), .config_in(config_chain[5697:5696])); 
mux4 mux_546 (.in({n2717, n1776, n1267, n1252}), .out(n1796), .config_in(config_chain[5699:5698])); 
mux3 mux_547 (.in({n2825, n1267, n1252}), .out(n1797), .config_in(config_chain[5701:5700])); 
mux4 mux_548 (.in({n2719, n1778, n1270, n1255}), .out(n1798), .config_in(config_chain[5703:5702])); 
mux3 mux_549 (.in({n2823, n1270, n1255}), .out(n1799), .config_in(config_chain[5705:5704])); 
mux4 mux_550 (.in({n2721, n1780, n1270, n1255}), .out(n1800), .config_in(config_chain[5707:5706])); 
mux3 mux_551 (.in({n2821, n1270, n1255}), .out(n1801), .config_in(config_chain[5709:5708])); 
mux3 mux_552 (.in({n2723, n1782, n1258}), .out(n1802), .config_in(config_chain[5711:5710])); 
mux2 mux_553 (.in({n2819, n1258}), .out(n1803), .config_in(config_chain[5712:5712])); 
mux3 mux_554 (.in({n2725, n1784, n1258}), .out(n1804), .config_in(config_chain[5714:5713])); 
mux2 mux_555 (.in({n2817, n1258}), .out(n1805), .config_in(config_chain[5715:5715])); 
mux3 mux_556 (.in({n2727, n1786, n1261}), .out(n1806), .config_in(config_chain[5717:5716])); 
mux2 mux_557 (.in({n2815, n1261}), .out(n1807), .config_in(config_chain[5718:5718])); 
mux3 mux_558 (.in({n2729, n1788, n1261}), .out(n1808), .config_in(config_chain[5720:5719])); 
mux2 mux_559 (.in({n2813, n1261}), .out(n1809), .config_in(config_chain[5721:5721])); 
mux3 mux_560 (.in({n2337, n2316, n315}), .out(n1810), .config_in(config_chain[5723:5722])); 
mux4 mux_561 (.in({n2431, n2428, n1831, n315}), .out(n1811), .config_in(config_chain[5725:5724])); 
mux3 mux_562 (.in({n2339, n2318, n315}), .out(n1812), .config_in(config_chain[5727:5726])); 
mux4 mux_563 (.in({n2449, n2410, n1833, n315}), .out(n1813), .config_in(config_chain[5729:5728])); 
mux2 mux_564 (.in({n2331, n2310}), .out(n1814), .config_in(config_chain[5730:5730])); 
mux3 mux_565 (.in({n2447, n2412, n1835}), .out(n1815), .config_in(config_chain[5732:5731])); 
mux2 mux_566 (.in({n2341, n2320}), .out(n1816), .config_in(config_chain[5733:5733])); 
mux3 mux_567 (.in({n2445, n2414, n1837}), .out(n1817), .config_in(config_chain[5735:5734])); 
mux2 mux_568 (.in({n2343, n2322}), .out(n1818), .config_in(config_chain[5736:5736])); 
mux3 mux_569 (.in({n2443, n2416, n1839}), .out(n1819), .config_in(config_chain[5738:5737])); 
mux2 mux_570 (.in({n2333, n2312}), .out(n1820), .config_in(config_chain[5739:5739])); 
mux3 mux_571 (.in({n2441, n2418, n1841}), .out(n1821), .config_in(config_chain[5741:5740])); 
mux2 mux_572 (.in({n2345, n2324}), .out(n1822), .config_in(config_chain[5742:5742])); 
mux3 mux_573 (.in({n2439, n2420, n1843}), .out(n1823), .config_in(config_chain[5744:5743])); 
mux2 mux_574 (.in({n2347, n2326}), .out(n1824), .config_in(config_chain[5745:5745])); 
mux3 mux_575 (.in({n2437, n2422, n1845}), .out(n1825), .config_in(config_chain[5747:5746])); 
mux2 mux_576 (.in({n2335, n2314}), .out(n1826), .config_in(config_chain[5748:5748])); 
mux3 mux_577 (.in({n2435, n2424, n1847}), .out(n1827), .config_in(config_chain[5750:5749])); 
mux2 mux_578 (.in({n2349, n2328}), .out(n1828), .config_in(config_chain[5751:5751])); 
mux3 mux_579 (.in({n2433, n2426, n1849}), .out(n1829), .config_in(config_chain[5753:5752])); 
mux4 mux_580 (.in({n2449, n2426, n1810, n561}), .out(n1830), .config_in(config_chain[5755:5754])); 
mux4 mux_581 (.in({n2531, n2528, n1851, n561}), .out(n1831), .config_in(config_chain[5757:5756])); 
mux4 mux_582 (.in({n2431, n2424, n1812, n561}), .out(n1832), .config_in(config_chain[5759:5758])); 
mux4 mux_583 (.in({n2549, n2510, n1853, n561}), .out(n1833), .config_in(config_chain[5761:5760])); 
mux3 mux_584 (.in({n2433, n2422, n1814}), .out(n1834), .config_in(config_chain[5763:5762])); 
mux3 mux_585 (.in({n2547, n2512, n1855}), .out(n1835), .config_in(config_chain[5765:5764])); 
mux3 mux_586 (.in({n2435, n2420, n1816}), .out(n1836), .config_in(config_chain[5767:5766])); 
mux3 mux_587 (.in({n2545, n2514, n1857}), .out(n1837), .config_in(config_chain[5769:5768])); 
mux3 mux_588 (.in({n2437, n2418, n1818}), .out(n1838), .config_in(config_chain[5771:5770])); 
mux3 mux_589 (.in({n2543, n2516, n1859}), .out(n1839), .config_in(config_chain[5773:5772])); 
mux3 mux_590 (.in({n2439, n2416, n1820}), .out(n1840), .config_in(config_chain[5775:5774])); 
mux3 mux_591 (.in({n2541, n2518, n1861}), .out(n1841), .config_in(config_chain[5777:5776])); 
mux3 mux_592 (.in({n2441, n2414, n1822}), .out(n1842), .config_in(config_chain[5779:5778])); 
mux3 mux_593 (.in({n2539, n2520, n1863}), .out(n1843), .config_in(config_chain[5781:5780])); 
mux3 mux_594 (.in({n2443, n2412, n1824}), .out(n1844), .config_in(config_chain[5783:5782])); 
mux3 mux_595 (.in({n2537, n2522, n1865}), .out(n1845), .config_in(config_chain[5785:5784])); 
mux3 mux_596 (.in({n2445, n2410, n1826}), .out(n1846), .config_in(config_chain[5787:5786])); 
mux3 mux_597 (.in({n2535, n2524, n1867}), .out(n1847), .config_in(config_chain[5789:5788])); 
mux3 mux_598 (.in({n2447, n2428, n1828}), .out(n1848), .config_in(config_chain[5791:5790])); 
mux3 mux_599 (.in({n2533, n2526, n1869}), .out(n1849), .config_in(config_chain[5793:5792])); 
mux4 mux_600 (.in({n2549, n2526, n1830, n807}), .out(n1850), .config_in(config_chain[5795:5794])); 
mux4 mux_601 (.in({n2631, n2628, n1871, n807}), .out(n1851), .config_in(config_chain[5797:5796])); 
mux4 mux_602 (.in({n2531, n2524, n1832, n807}), .out(n1852), .config_in(config_chain[5799:5798])); 
mux4 mux_603 (.in({n2649, n2610, n1873, n807}), .out(n1853), .config_in(config_chain[5801:5800])); 
mux3 mux_604 (.in({n2533, n2522, n1834}), .out(n1854), .config_in(config_chain[5803:5802])); 
mux3 mux_605 (.in({n2647, n2612, n1875}), .out(n1855), .config_in(config_chain[5805:5804])); 
mux3 mux_606 (.in({n2535, n2520, n1836}), .out(n1856), .config_in(config_chain[5807:5806])); 
mux3 mux_607 (.in({n2645, n2614, n1877}), .out(n1857), .config_in(config_chain[5809:5808])); 
mux3 mux_608 (.in({n2537, n2518, n1838}), .out(n1858), .config_in(config_chain[5811:5810])); 
mux3 mux_609 (.in({n2643, n2616, n1879}), .out(n1859), .config_in(config_chain[5813:5812])); 
mux3 mux_610 (.in({n2539, n2516, n1840}), .out(n1860), .config_in(config_chain[5815:5814])); 
mux3 mux_611 (.in({n2641, n2618, n1881}), .out(n1861), .config_in(config_chain[5817:5816])); 
mux3 mux_612 (.in({n2541, n2514, n1842}), .out(n1862), .config_in(config_chain[5819:5818])); 
mux3 mux_613 (.in({n2639, n2620, n1883}), .out(n1863), .config_in(config_chain[5821:5820])); 
mux3 mux_614 (.in({n2543, n2512, n1844}), .out(n1864), .config_in(config_chain[5823:5822])); 
mux3 mux_615 (.in({n2637, n2622, n1885}), .out(n1865), .config_in(config_chain[5825:5824])); 
mux3 mux_616 (.in({n2545, n2510, n1846}), .out(n1866), .config_in(config_chain[5827:5826])); 
mux3 mux_617 (.in({n2635, n2624, n1887}), .out(n1867), .config_in(config_chain[5829:5828])); 
mux3 mux_618 (.in({n2547, n2528, n1848}), .out(n1868), .config_in(config_chain[5831:5830])); 
mux3 mux_619 (.in({n2633, n2626, n1889}), .out(n1869), .config_in(config_chain[5833:5832])); 
mux4 mux_620 (.in({n2649, n2626, n1850, n1053}), .out(n1870), .config_in(config_chain[5835:5834])); 
mux4 mux_621 (.in({n2731, n2728, n1891, n1053}), .out(n1871), .config_in(config_chain[5837:5836])); 
mux4 mux_622 (.in({n2631, n2624, n1852, n1053}), .out(n1872), .config_in(config_chain[5839:5838])); 
mux4 mux_623 (.in({n2749, n2710, n1893, n1053}), .out(n1873), .config_in(config_chain[5841:5840])); 
mux3 mux_624 (.in({n2633, n2622, n1854}), .out(n1874), .config_in(config_chain[5843:5842])); 
mux3 mux_625 (.in({n2747, n2712, n1895}), .out(n1875), .config_in(config_chain[5845:5844])); 
mux3 mux_626 (.in({n2635, n2620, n1856}), .out(n1876), .config_in(config_chain[5847:5846])); 
mux3 mux_627 (.in({n2745, n2714, n1897}), .out(n1877), .config_in(config_chain[5849:5848])); 
mux3 mux_628 (.in({n2637, n2618, n1858}), .out(n1878), .config_in(config_chain[5851:5850])); 
mux3 mux_629 (.in({n2743, n2716, n1899}), .out(n1879), .config_in(config_chain[5853:5852])); 
mux3 mux_630 (.in({n2639, n2616, n1860}), .out(n1880), .config_in(config_chain[5855:5854])); 
mux3 mux_631 (.in({n2741, n2718, n1901}), .out(n1881), .config_in(config_chain[5857:5856])); 
mux3 mux_632 (.in({n2641, n2614, n1862}), .out(n1882), .config_in(config_chain[5859:5858])); 
mux3 mux_633 (.in({n2739, n2720, n1903}), .out(n1883), .config_in(config_chain[5861:5860])); 
mux3 mux_634 (.in({n2643, n2612, n1864}), .out(n1884), .config_in(config_chain[5863:5862])); 
mux3 mux_635 (.in({n2737, n2722, n1905}), .out(n1885), .config_in(config_chain[5865:5864])); 
mux3 mux_636 (.in({n2645, n2610, n1866}), .out(n1886), .config_in(config_chain[5867:5866])); 
mux3 mux_637 (.in({n2735, n2724, n1907}), .out(n1887), .config_in(config_chain[5869:5868])); 
mux3 mux_638 (.in({n2647, n2628, n1868}), .out(n1888), .config_in(config_chain[5871:5870])); 
mux3 mux_639 (.in({n2733, n2726, n1909}), .out(n1889), .config_in(config_chain[5873:5872])); 
mux4 mux_640 (.in({n2749, n2726, n1870, n1299}), .out(n1890), .config_in(config_chain[5875:5874])); 
mux3 mux_641 (.in({n2831, n2810, n1299}), .out(n1891), .config_in(config_chain[5877:5876])); 
mux4 mux_642 (.in({n2731, n2724, n1872, n1299}), .out(n1892), .config_in(config_chain[5879:5878])); 
mux3 mux_643 (.in({n2839, n2818, n1299}), .out(n1893), .config_in(config_chain[5881:5880])); 
mux3 mux_644 (.in({n2733, n2722, n1874}), .out(n1894), .config_in(config_chain[5883:5882])); 
mux2 mux_645 (.in({n2841, n2820}), .out(n1895), .config_in(config_chain[5884:5884])); 
mux3 mux_646 (.in({n2735, n2720, n1876}), .out(n1896), .config_in(config_chain[5886:5885])); 
mux2 mux_647 (.in({n2833, n2812}), .out(n1897), .config_in(config_chain[5887:5887])); 
mux3 mux_648 (.in({n2737, n2718, n1878}), .out(n1898), .config_in(config_chain[5889:5888])); 
mux2 mux_649 (.in({n2843, n2822}), .out(n1899), .config_in(config_chain[5890:5890])); 
mux3 mux_650 (.in({n2739, n2716, n1880}), .out(n1900), .config_in(config_chain[5892:5891])); 
mux2 mux_651 (.in({n2845, n2824}), .out(n1901), .config_in(config_chain[5893:5893])); 
mux3 mux_652 (.in({n2741, n2714, n1882}), .out(n1902), .config_in(config_chain[5895:5894])); 
mux2 mux_653 (.in({n2835, n2814}), .out(n1903), .config_in(config_chain[5896:5896])); 
mux3 mux_654 (.in({n2743, n2712, n1884}), .out(n1904), .config_in(config_chain[5898:5897])); 
mux2 mux_655 (.in({n2847, n2826}), .out(n1905), .config_in(config_chain[5899:5899])); 
mux3 mux_656 (.in({n2745, n2710, n1886}), .out(n1906), .config_in(config_chain[5901:5900])); 
mux2 mux_657 (.in({n2849, n2828}), .out(n1907), .config_in(config_chain[5902:5902])); 
mux3 mux_658 (.in({n2747, n2728, n1888}), .out(n1908), .config_in(config_chain[5904:5903])); 
mux2 mux_659 (.in({n2837, n2816}), .out(n1909), .config_in(config_chain[5905:5905])); 
mux3 mux_660 (.in({n2357, n2336, n345}), .out(n1910), .config_in(config_chain[5907:5906])); 
mux4 mux_661 (.in({n2451, n2448, n1931, n345}), .out(n1911), .config_in(config_chain[5909:5908])); 
mux3 mux_662 (.in({n2359, n2338, n345}), .out(n1912), .config_in(config_chain[5911:5910])); 
mux4 mux_663 (.in({n2469, n2430, n1933, n345}), .out(n1913), .config_in(config_chain[5913:5912])); 
mux2 mux_664 (.in({n2351, n2330}), .out(n1914), .config_in(config_chain[5914:5914])); 
mux3 mux_665 (.in({n2467, n2432, n1935}), .out(n1915), .config_in(config_chain[5916:5915])); 
mux2 mux_666 (.in({n2361, n2340}), .out(n1916), .config_in(config_chain[5917:5917])); 
mux3 mux_667 (.in({n2465, n2434, n1937}), .out(n1917), .config_in(config_chain[5919:5918])); 
mux2 mux_668 (.in({n2363, n2342}), .out(n1918), .config_in(config_chain[5920:5920])); 
mux3 mux_669 (.in({n2463, n2436, n1939}), .out(n1919), .config_in(config_chain[5922:5921])); 
mux2 mux_670 (.in({n2353, n2332}), .out(n1920), .config_in(config_chain[5923:5923])); 
mux3 mux_671 (.in({n2461, n2438, n1941}), .out(n1921), .config_in(config_chain[5925:5924])); 
mux2 mux_672 (.in({n2365, n2344}), .out(n1922), .config_in(config_chain[5926:5926])); 
mux3 mux_673 (.in({n2459, n2440, n1943}), .out(n1923), .config_in(config_chain[5928:5927])); 
mux2 mux_674 (.in({n2367, n2346}), .out(n1924), .config_in(config_chain[5929:5929])); 
mux3 mux_675 (.in({n2457, n2442, n1945}), .out(n1925), .config_in(config_chain[5931:5930])); 
mux2 mux_676 (.in({n2355, n2334}), .out(n1926), .config_in(config_chain[5932:5932])); 
mux3 mux_677 (.in({n2455, n2444, n1947}), .out(n1927), .config_in(config_chain[5934:5933])); 
mux2 mux_678 (.in({n2369, n2348}), .out(n1928), .config_in(config_chain[5935:5935])); 
mux3 mux_679 (.in({n2453, n2446, n1949}), .out(n1929), .config_in(config_chain[5937:5936])); 
mux4 mux_680 (.in({n2469, n2446, n1910, n591}), .out(n1930), .config_in(config_chain[5939:5938])); 
mux4 mux_681 (.in({n2551, n2548, n1951, n591}), .out(n1931), .config_in(config_chain[5941:5940])); 
mux4 mux_682 (.in({n2451, n2444, n1912, n591}), .out(n1932), .config_in(config_chain[5943:5942])); 
mux4 mux_683 (.in({n2569, n2530, n1953, n591}), .out(n1933), .config_in(config_chain[5945:5944])); 
mux3 mux_684 (.in({n2453, n2442, n1914}), .out(n1934), .config_in(config_chain[5947:5946])); 
mux3 mux_685 (.in({n2567, n2532, n1955}), .out(n1935), .config_in(config_chain[5949:5948])); 
mux3 mux_686 (.in({n2455, n2440, n1916}), .out(n1936), .config_in(config_chain[5951:5950])); 
mux3 mux_687 (.in({n2565, n2534, n1957}), .out(n1937), .config_in(config_chain[5953:5952])); 
mux3 mux_688 (.in({n2457, n2438, n1918}), .out(n1938), .config_in(config_chain[5955:5954])); 
mux3 mux_689 (.in({n2563, n2536, n1959}), .out(n1939), .config_in(config_chain[5957:5956])); 
mux3 mux_690 (.in({n2459, n2436, n1920}), .out(n1940), .config_in(config_chain[5959:5958])); 
mux3 mux_691 (.in({n2561, n2538, n1961}), .out(n1941), .config_in(config_chain[5961:5960])); 
mux3 mux_692 (.in({n2461, n2434, n1922}), .out(n1942), .config_in(config_chain[5963:5962])); 
mux3 mux_693 (.in({n2559, n2540, n1963}), .out(n1943), .config_in(config_chain[5965:5964])); 
mux3 mux_694 (.in({n2463, n2432, n1924}), .out(n1944), .config_in(config_chain[5967:5966])); 
mux3 mux_695 (.in({n2557, n2542, n1965}), .out(n1945), .config_in(config_chain[5969:5968])); 
mux3 mux_696 (.in({n2465, n2430, n1926}), .out(n1946), .config_in(config_chain[5971:5970])); 
mux3 mux_697 (.in({n2555, n2544, n1967}), .out(n1947), .config_in(config_chain[5973:5972])); 
mux3 mux_698 (.in({n2467, n2448, n1928}), .out(n1948), .config_in(config_chain[5975:5974])); 
mux3 mux_699 (.in({n2553, n2546, n1969}), .out(n1949), .config_in(config_chain[5977:5976])); 
mux4 mux_700 (.in({n2569, n2546, n1930, n837}), .out(n1950), .config_in(config_chain[5979:5978])); 
mux4 mux_701 (.in({n2651, n2648, n1971, n837}), .out(n1951), .config_in(config_chain[5981:5980])); 
mux4 mux_702 (.in({n2551, n2544, n1932, n837}), .out(n1952), .config_in(config_chain[5983:5982])); 
mux4 mux_703 (.in({n2669, n2630, n1973, n837}), .out(n1953), .config_in(config_chain[5985:5984])); 
mux3 mux_704 (.in({n2553, n2542, n1934}), .out(n1954), .config_in(config_chain[5987:5986])); 
mux3 mux_705 (.in({n2667, n2632, n1975}), .out(n1955), .config_in(config_chain[5989:5988])); 
mux3 mux_706 (.in({n2555, n2540, n1936}), .out(n1956), .config_in(config_chain[5991:5990])); 
mux3 mux_707 (.in({n2665, n2634, n1977}), .out(n1957), .config_in(config_chain[5993:5992])); 
mux3 mux_708 (.in({n2557, n2538, n1938}), .out(n1958), .config_in(config_chain[5995:5994])); 
mux3 mux_709 (.in({n2663, n2636, n1979}), .out(n1959), .config_in(config_chain[5997:5996])); 
mux3 mux_710 (.in({n2559, n2536, n1940}), .out(n1960), .config_in(config_chain[5999:5998])); 
mux3 mux_711 (.in({n2661, n2638, n1981}), .out(n1961), .config_in(config_chain[6001:6000])); 
mux3 mux_712 (.in({n2561, n2534, n1942}), .out(n1962), .config_in(config_chain[6003:6002])); 
mux3 mux_713 (.in({n2659, n2640, n1983}), .out(n1963), .config_in(config_chain[6005:6004])); 
mux3 mux_714 (.in({n2563, n2532, n1944}), .out(n1964), .config_in(config_chain[6007:6006])); 
mux3 mux_715 (.in({n2657, n2642, n1985}), .out(n1965), .config_in(config_chain[6009:6008])); 
mux3 mux_716 (.in({n2565, n2530, n1946}), .out(n1966), .config_in(config_chain[6011:6010])); 
mux3 mux_717 (.in({n2655, n2644, n1987}), .out(n1967), .config_in(config_chain[6013:6012])); 
mux3 mux_718 (.in({n2567, n2548, n1948}), .out(n1968), .config_in(config_chain[6015:6014])); 
mux3 mux_719 (.in({n2653, n2646, n1989}), .out(n1969), .config_in(config_chain[6017:6016])); 
mux4 mux_720 (.in({n2669, n2646, n1950, n1083}), .out(n1970), .config_in(config_chain[6019:6018])); 
mux4 mux_721 (.in({n2751, n2748, n1991, n1083}), .out(n1971), .config_in(config_chain[6021:6020])); 
mux4 mux_722 (.in({n2651, n2644, n1952, n1083}), .out(n1972), .config_in(config_chain[6023:6022])); 
mux4 mux_723 (.in({n2769, n2730, n1993, n1083}), .out(n1973), .config_in(config_chain[6025:6024])); 
mux3 mux_724 (.in({n2653, n2642, n1954}), .out(n1974), .config_in(config_chain[6027:6026])); 
mux3 mux_725 (.in({n2767, n2732, n1995}), .out(n1975), .config_in(config_chain[6029:6028])); 
mux3 mux_726 (.in({n2655, n2640, n1956}), .out(n1976), .config_in(config_chain[6031:6030])); 
mux3 mux_727 (.in({n2765, n2734, n1997}), .out(n1977), .config_in(config_chain[6033:6032])); 
mux3 mux_728 (.in({n2657, n2638, n1958}), .out(n1978), .config_in(config_chain[6035:6034])); 
mux3 mux_729 (.in({n2763, n2736, n1999}), .out(n1979), .config_in(config_chain[6037:6036])); 
mux3 mux_730 (.in({n2659, n2636, n1960}), .out(n1980), .config_in(config_chain[6039:6038])); 
mux3 mux_731 (.in({n2761, n2738, n2001}), .out(n1981), .config_in(config_chain[6041:6040])); 
mux3 mux_732 (.in({n2661, n2634, n1962}), .out(n1982), .config_in(config_chain[6043:6042])); 
mux3 mux_733 (.in({n2759, n2740, n2003}), .out(n1983), .config_in(config_chain[6045:6044])); 
mux3 mux_734 (.in({n2663, n2632, n1964}), .out(n1984), .config_in(config_chain[6047:6046])); 
mux3 mux_735 (.in({n2757, n2742, n2005}), .out(n1985), .config_in(config_chain[6049:6048])); 
mux3 mux_736 (.in({n2665, n2630, n1966}), .out(n1986), .config_in(config_chain[6051:6050])); 
mux3 mux_737 (.in({n2755, n2744, n2007}), .out(n1987), .config_in(config_chain[6053:6052])); 
mux3 mux_738 (.in({n2667, n2648, n1968}), .out(n1988), .config_in(config_chain[6055:6054])); 
mux3 mux_739 (.in({n2753, n2746, n2009}), .out(n1989), .config_in(config_chain[6057:6056])); 
mux4 mux_740 (.in({n2769, n2746, n1970, n1329}), .out(n1990), .config_in(config_chain[6059:6058])); 
mux3 mux_741 (.in({n2851, n2830, n1329}), .out(n1991), .config_in(config_chain[6061:6060])); 
mux4 mux_742 (.in({n2751, n2744, n1972, n1329}), .out(n1992), .config_in(config_chain[6063:6062])); 
mux3 mux_743 (.in({n2859, n2838, n1329}), .out(n1993), .config_in(config_chain[6065:6064])); 
mux3 mux_744 (.in({n2753, n2742, n1974}), .out(n1994), .config_in(config_chain[6067:6066])); 
mux2 mux_745 (.in({n2861, n2840}), .out(n1995), .config_in(config_chain[6068:6068])); 
mux3 mux_746 (.in({n2755, n2740, n1976}), .out(n1996), .config_in(config_chain[6070:6069])); 
mux2 mux_747 (.in({n2853, n2832}), .out(n1997), .config_in(config_chain[6071:6071])); 
mux3 mux_748 (.in({n2757, n2738, n1978}), .out(n1998), .config_in(config_chain[6073:6072])); 
mux2 mux_749 (.in({n2863, n2842}), .out(n1999), .config_in(config_chain[6074:6074])); 
mux3 mux_750 (.in({n2759, n2736, n1980}), .out(n2000), .config_in(config_chain[6076:6075])); 
mux2 mux_751 (.in({n2865, n2844}), .out(n2001), .config_in(config_chain[6077:6077])); 
mux3 mux_752 (.in({n2761, n2734, n1982}), .out(n2002), .config_in(config_chain[6079:6078])); 
mux2 mux_753 (.in({n2855, n2834}), .out(n2003), .config_in(config_chain[6080:6080])); 
mux3 mux_754 (.in({n2763, n2732, n1984}), .out(n2004), .config_in(config_chain[6082:6081])); 
mux2 mux_755 (.in({n2867, n2846}), .out(n2005), .config_in(config_chain[6083:6083])); 
mux3 mux_756 (.in({n2765, n2730, n1986}), .out(n2006), .config_in(config_chain[6085:6084])); 
mux2 mux_757 (.in({n2869, n2848}), .out(n2007), .config_in(config_chain[6086:6086])); 
mux3 mux_758 (.in({n2767, n2748, n1988}), .out(n2008), .config_in(config_chain[6088:6087])); 
mux2 mux_759 (.in({n2857, n2836}), .out(n2009), .config_in(config_chain[6089:6089])); 
mux3 mux_760 (.in({n2377, n2356, n375}), .out(n2010), .config_in(config_chain[6091:6090])); 
mux4 mux_761 (.in({n2471, n2468, n2031, n375}), .out(n2011), .config_in(config_chain[6093:6092])); 
mux3 mux_762 (.in({n2379, n2358, n375}), .out(n2012), .config_in(config_chain[6095:6094])); 
mux4 mux_763 (.in({n2489, n2450, n2033, n375}), .out(n2013), .config_in(config_chain[6097:6096])); 
mux2 mux_764 (.in({n2371, n2350}), .out(n2014), .config_in(config_chain[6098:6098])); 
mux3 mux_765 (.in({n2487, n2452, n2035}), .out(n2015), .config_in(config_chain[6100:6099])); 
mux2 mux_766 (.in({n2381, n2360}), .out(n2016), .config_in(config_chain[6101:6101])); 
mux3 mux_767 (.in({n2485, n2454, n2037}), .out(n2017), .config_in(config_chain[6103:6102])); 
mux2 mux_768 (.in({n2383, n2362}), .out(n2018), .config_in(config_chain[6104:6104])); 
mux3 mux_769 (.in({n2483, n2456, n2039}), .out(n2019), .config_in(config_chain[6106:6105])); 
mux2 mux_770 (.in({n2373, n2352}), .out(n2020), .config_in(config_chain[6107:6107])); 
mux3 mux_771 (.in({n2481, n2458, n2041}), .out(n2021), .config_in(config_chain[6109:6108])); 
mux2 mux_772 (.in({n2385, n2364}), .out(n2022), .config_in(config_chain[6110:6110])); 
mux3 mux_773 (.in({n2479, n2460, n2043}), .out(n2023), .config_in(config_chain[6112:6111])); 
mux2 mux_774 (.in({n2387, n2366}), .out(n2024), .config_in(config_chain[6113:6113])); 
mux3 mux_775 (.in({n2477, n2462, n2045}), .out(n2025), .config_in(config_chain[6115:6114])); 
mux2 mux_776 (.in({n2375, n2354}), .out(n2026), .config_in(config_chain[6116:6116])); 
mux3 mux_777 (.in({n2475, n2464, n2047}), .out(n2027), .config_in(config_chain[6118:6117])); 
mux2 mux_778 (.in({n2389, n2368}), .out(n2028), .config_in(config_chain[6119:6119])); 
mux3 mux_779 (.in({n2473, n2466, n2049}), .out(n2029), .config_in(config_chain[6121:6120])); 
mux4 mux_780 (.in({n2489, n2466, n2010, n621}), .out(n2030), .config_in(config_chain[6123:6122])); 
mux4 mux_781 (.in({n2571, n2568, n2051, n621}), .out(n2031), .config_in(config_chain[6125:6124])); 
mux4 mux_782 (.in({n2471, n2464, n2012, n621}), .out(n2032), .config_in(config_chain[6127:6126])); 
mux4 mux_783 (.in({n2589, n2550, n2053, n621}), .out(n2033), .config_in(config_chain[6129:6128])); 
mux3 mux_784 (.in({n2473, n2462, n2014}), .out(n2034), .config_in(config_chain[6131:6130])); 
mux3 mux_785 (.in({n2587, n2552, n2055}), .out(n2035), .config_in(config_chain[6133:6132])); 
mux3 mux_786 (.in({n2475, n2460, n2016}), .out(n2036), .config_in(config_chain[6135:6134])); 
mux3 mux_787 (.in({n2585, n2554, n2057}), .out(n2037), .config_in(config_chain[6137:6136])); 
mux3 mux_788 (.in({n2477, n2458, n2018}), .out(n2038), .config_in(config_chain[6139:6138])); 
mux3 mux_789 (.in({n2583, n2556, n2059}), .out(n2039), .config_in(config_chain[6141:6140])); 
mux3 mux_790 (.in({n2479, n2456, n2020}), .out(n2040), .config_in(config_chain[6143:6142])); 
mux3 mux_791 (.in({n2581, n2558, n2061}), .out(n2041), .config_in(config_chain[6145:6144])); 
mux3 mux_792 (.in({n2481, n2454, n2022}), .out(n2042), .config_in(config_chain[6147:6146])); 
mux3 mux_793 (.in({n2579, n2560, n2063}), .out(n2043), .config_in(config_chain[6149:6148])); 
mux3 mux_794 (.in({n2483, n2452, n2024}), .out(n2044), .config_in(config_chain[6151:6150])); 
mux3 mux_795 (.in({n2577, n2562, n2065}), .out(n2045), .config_in(config_chain[6153:6152])); 
mux3 mux_796 (.in({n2485, n2450, n2026}), .out(n2046), .config_in(config_chain[6155:6154])); 
mux3 mux_797 (.in({n2575, n2564, n2067}), .out(n2047), .config_in(config_chain[6157:6156])); 
mux3 mux_798 (.in({n2487, n2468, n2028}), .out(n2048), .config_in(config_chain[6159:6158])); 
mux3 mux_799 (.in({n2573, n2566, n2069}), .out(n2049), .config_in(config_chain[6161:6160])); 
mux4 mux_800 (.in({n2589, n2566, n2030, n867}), .out(n2050), .config_in(config_chain[6163:6162])); 
mux4 mux_801 (.in({n2671, n2668, n2071, n867}), .out(n2051), .config_in(config_chain[6165:6164])); 
mux4 mux_802 (.in({n2571, n2564, n2032, n867}), .out(n2052), .config_in(config_chain[6167:6166])); 
mux4 mux_803 (.in({n2689, n2650, n2073, n867}), .out(n2053), .config_in(config_chain[6169:6168])); 
mux3 mux_804 (.in({n2573, n2562, n2034}), .out(n2054), .config_in(config_chain[6171:6170])); 
mux3 mux_805 (.in({n2687, n2652, n2075}), .out(n2055), .config_in(config_chain[6173:6172])); 
mux3 mux_806 (.in({n2575, n2560, n2036}), .out(n2056), .config_in(config_chain[6175:6174])); 
mux3 mux_807 (.in({n2685, n2654, n2077}), .out(n2057), .config_in(config_chain[6177:6176])); 
mux3 mux_808 (.in({n2577, n2558, n2038}), .out(n2058), .config_in(config_chain[6179:6178])); 
mux3 mux_809 (.in({n2683, n2656, n2079}), .out(n2059), .config_in(config_chain[6181:6180])); 
mux3 mux_810 (.in({n2579, n2556, n2040}), .out(n2060), .config_in(config_chain[6183:6182])); 
mux3 mux_811 (.in({n2681, n2658, n2081}), .out(n2061), .config_in(config_chain[6185:6184])); 
mux3 mux_812 (.in({n2581, n2554, n2042}), .out(n2062), .config_in(config_chain[6187:6186])); 
mux3 mux_813 (.in({n2679, n2660, n2083}), .out(n2063), .config_in(config_chain[6189:6188])); 
mux3 mux_814 (.in({n2583, n2552, n2044}), .out(n2064), .config_in(config_chain[6191:6190])); 
mux3 mux_815 (.in({n2677, n2662, n2085}), .out(n2065), .config_in(config_chain[6193:6192])); 
mux3 mux_816 (.in({n2585, n2550, n2046}), .out(n2066), .config_in(config_chain[6195:6194])); 
mux3 mux_817 (.in({n2675, n2664, n2087}), .out(n2067), .config_in(config_chain[6197:6196])); 
mux3 mux_818 (.in({n2587, n2568, n2048}), .out(n2068), .config_in(config_chain[6199:6198])); 
mux3 mux_819 (.in({n2673, n2666, n2089}), .out(n2069), .config_in(config_chain[6201:6200])); 
mux4 mux_820 (.in({n2689, n2666, n2050, n1113}), .out(n2070), .config_in(config_chain[6203:6202])); 
mux4 mux_821 (.in({n2771, n2768, n2091, n1113}), .out(n2071), .config_in(config_chain[6205:6204])); 
mux4 mux_822 (.in({n2671, n2664, n2052, n1113}), .out(n2072), .config_in(config_chain[6207:6206])); 
mux4 mux_823 (.in({n2789, n2750, n2093, n1113}), .out(n2073), .config_in(config_chain[6209:6208])); 
mux3 mux_824 (.in({n2673, n2662, n2054}), .out(n2074), .config_in(config_chain[6211:6210])); 
mux3 mux_825 (.in({n2787, n2752, n2095}), .out(n2075), .config_in(config_chain[6213:6212])); 
mux3 mux_826 (.in({n2675, n2660, n2056}), .out(n2076), .config_in(config_chain[6215:6214])); 
mux3 mux_827 (.in({n2785, n2754, n2097}), .out(n2077), .config_in(config_chain[6217:6216])); 
mux3 mux_828 (.in({n2677, n2658, n2058}), .out(n2078), .config_in(config_chain[6219:6218])); 
mux3 mux_829 (.in({n2783, n2756, n2099}), .out(n2079), .config_in(config_chain[6221:6220])); 
mux3 mux_830 (.in({n2679, n2656, n2060}), .out(n2080), .config_in(config_chain[6223:6222])); 
mux3 mux_831 (.in({n2781, n2758, n2101}), .out(n2081), .config_in(config_chain[6225:6224])); 
mux3 mux_832 (.in({n2681, n2654, n2062}), .out(n2082), .config_in(config_chain[6227:6226])); 
mux3 mux_833 (.in({n2779, n2760, n2103}), .out(n2083), .config_in(config_chain[6229:6228])); 
mux3 mux_834 (.in({n2683, n2652, n2064}), .out(n2084), .config_in(config_chain[6231:6230])); 
mux3 mux_835 (.in({n2777, n2762, n2105}), .out(n2085), .config_in(config_chain[6233:6232])); 
mux3 mux_836 (.in({n2685, n2650, n2066}), .out(n2086), .config_in(config_chain[6235:6234])); 
mux3 mux_837 (.in({n2775, n2764, n2107}), .out(n2087), .config_in(config_chain[6237:6236])); 
mux3 mux_838 (.in({n2687, n2668, n2068}), .out(n2088), .config_in(config_chain[6239:6238])); 
mux3 mux_839 (.in({n2773, n2766, n2109}), .out(n2089), .config_in(config_chain[6241:6240])); 
mux4 mux_840 (.in({n2789, n2766, n2070, n1359}), .out(n2090), .config_in(config_chain[6243:6242])); 
mux3 mux_841 (.in({n2871, n2850, n1359}), .out(n2091), .config_in(config_chain[6245:6244])); 
mux4 mux_842 (.in({n2771, n2764, n2072, n1359}), .out(n2092), .config_in(config_chain[6247:6246])); 
mux3 mux_843 (.in({n2879, n2858, n1359}), .out(n2093), .config_in(config_chain[6249:6248])); 
mux3 mux_844 (.in({n2773, n2762, n2074}), .out(n2094), .config_in(config_chain[6251:6250])); 
mux2 mux_845 (.in({n2881, n2860}), .out(n2095), .config_in(config_chain[6252:6252])); 
mux3 mux_846 (.in({n2775, n2760, n2076}), .out(n2096), .config_in(config_chain[6254:6253])); 
mux2 mux_847 (.in({n2873, n2852}), .out(n2097), .config_in(config_chain[6255:6255])); 
mux3 mux_848 (.in({n2777, n2758, n2078}), .out(n2098), .config_in(config_chain[6257:6256])); 
mux2 mux_849 (.in({n2883, n2862}), .out(n2099), .config_in(config_chain[6258:6258])); 
mux3 mux_850 (.in({n2779, n2756, n2080}), .out(n2100), .config_in(config_chain[6260:6259])); 
mux2 mux_851 (.in({n2885, n2864}), .out(n2101), .config_in(config_chain[6261:6261])); 
mux3 mux_852 (.in({n2781, n2754, n2082}), .out(n2102), .config_in(config_chain[6263:6262])); 
mux2 mux_853 (.in({n2875, n2854}), .out(n2103), .config_in(config_chain[6264:6264])); 
mux3 mux_854 (.in({n2783, n2752, n2084}), .out(n2104), .config_in(config_chain[6266:6265])); 
mux2 mux_855 (.in({n2887, n2866}), .out(n2105), .config_in(config_chain[6267:6267])); 
mux3 mux_856 (.in({n2785, n2750, n2086}), .out(n2106), .config_in(config_chain[6269:6268])); 
mux2 mux_857 (.in({n2889, n2868}), .out(n2107), .config_in(config_chain[6270:6270])); 
mux3 mux_858 (.in({n2787, n2768, n2088}), .out(n2108), .config_in(config_chain[6272:6271])); 
mux2 mux_859 (.in({n2877, n2856}), .out(n2109), .config_in(config_chain[6273:6273])); 
mux3 mux_860 (.in({n2397, n2376, n405}), .out(n2110), .config_in(config_chain[6275:6274])); 
mux4 mux_861 (.in({n2491, n2488, n2131, n405}), .out(n2111), .config_in(config_chain[6277:6276])); 
mux3 mux_862 (.in({n2399, n2378, n405}), .out(n2112), .config_in(config_chain[6279:6278])); 
mux4 mux_863 (.in({n2509, n2470, n2133, n405}), .out(n2113), .config_in(config_chain[6281:6280])); 
mux2 mux_864 (.in({n2391, n2370}), .out(n2114), .config_in(config_chain[6282:6282])); 
mux3 mux_865 (.in({n2507, n2472, n2135}), .out(n2115), .config_in(config_chain[6284:6283])); 
mux2 mux_866 (.in({n2401, n2380}), .out(n2116), .config_in(config_chain[6285:6285])); 
mux3 mux_867 (.in({n2505, n2474, n2137}), .out(n2117), .config_in(config_chain[6287:6286])); 
mux2 mux_868 (.in({n2403, n2382}), .out(n2118), .config_in(config_chain[6288:6288])); 
mux3 mux_869 (.in({n2503, n2476, n2139}), .out(n2119), .config_in(config_chain[6290:6289])); 
mux2 mux_870 (.in({n2393, n2372}), .out(n2120), .config_in(config_chain[6291:6291])); 
mux3 mux_871 (.in({n2501, n2478, n2141}), .out(n2121), .config_in(config_chain[6293:6292])); 
mux2 mux_872 (.in({n2405, n2384}), .out(n2122), .config_in(config_chain[6294:6294])); 
mux3 mux_873 (.in({n2499, n2480, n2143}), .out(n2123), .config_in(config_chain[6296:6295])); 
mux2 mux_874 (.in({n2407, n2386}), .out(n2124), .config_in(config_chain[6297:6297])); 
mux3 mux_875 (.in({n2497, n2482, n2145}), .out(n2125), .config_in(config_chain[6299:6298])); 
mux2 mux_876 (.in({n2395, n2374}), .out(n2126), .config_in(config_chain[6300:6300])); 
mux3 mux_877 (.in({n2495, n2484, n2147}), .out(n2127), .config_in(config_chain[6302:6301])); 
mux2 mux_878 (.in({n2409, n2388}), .out(n2128), .config_in(config_chain[6303:6303])); 
mux3 mux_879 (.in({n2493, n2486, n2149}), .out(n2129), .config_in(config_chain[6305:6304])); 
mux4 mux_880 (.in({n2509, n2486, n2110, n651}), .out(n2130), .config_in(config_chain[6307:6306])); 
mux4 mux_881 (.in({n2591, n2588, n2151, n651}), .out(n2131), .config_in(config_chain[6309:6308])); 
mux4 mux_882 (.in({n2491, n2484, n2112, n651}), .out(n2132), .config_in(config_chain[6311:6310])); 
mux4 mux_883 (.in({n2609, n2570, n2153, n651}), .out(n2133), .config_in(config_chain[6313:6312])); 
mux3 mux_884 (.in({n2493, n2482, n2114}), .out(n2134), .config_in(config_chain[6315:6314])); 
mux3 mux_885 (.in({n2607, n2572, n2155}), .out(n2135), .config_in(config_chain[6317:6316])); 
mux3 mux_886 (.in({n2495, n2480, n2116}), .out(n2136), .config_in(config_chain[6319:6318])); 
mux3 mux_887 (.in({n2605, n2574, n2157}), .out(n2137), .config_in(config_chain[6321:6320])); 
mux3 mux_888 (.in({n2497, n2478, n2118}), .out(n2138), .config_in(config_chain[6323:6322])); 
mux3 mux_889 (.in({n2603, n2576, n2159}), .out(n2139), .config_in(config_chain[6325:6324])); 
mux3 mux_890 (.in({n2499, n2476, n2120}), .out(n2140), .config_in(config_chain[6327:6326])); 
mux3 mux_891 (.in({n2601, n2578, n2161}), .out(n2141), .config_in(config_chain[6329:6328])); 
mux3 mux_892 (.in({n2501, n2474, n2122}), .out(n2142), .config_in(config_chain[6331:6330])); 
mux3 mux_893 (.in({n2599, n2580, n2163}), .out(n2143), .config_in(config_chain[6333:6332])); 
mux3 mux_894 (.in({n2503, n2472, n2124}), .out(n2144), .config_in(config_chain[6335:6334])); 
mux3 mux_895 (.in({n2597, n2582, n2165}), .out(n2145), .config_in(config_chain[6337:6336])); 
mux3 mux_896 (.in({n2505, n2470, n2126}), .out(n2146), .config_in(config_chain[6339:6338])); 
mux3 mux_897 (.in({n2595, n2584, n2167}), .out(n2147), .config_in(config_chain[6341:6340])); 
mux3 mux_898 (.in({n2507, n2488, n2128}), .out(n2148), .config_in(config_chain[6343:6342])); 
mux3 mux_899 (.in({n2593, n2586, n2169}), .out(n2149), .config_in(config_chain[6345:6344])); 
mux4 mux_900 (.in({n2609, n2586, n2130, n897}), .out(n2150), .config_in(config_chain[6347:6346])); 
mux4 mux_901 (.in({n2691, n2688, n2171, n897}), .out(n2151), .config_in(config_chain[6349:6348])); 
mux4 mux_902 (.in({n2591, n2584, n2132, n897}), .out(n2152), .config_in(config_chain[6351:6350])); 
mux4 mux_903 (.in({n2709, n2670, n2173, n897}), .out(n2153), .config_in(config_chain[6353:6352])); 
mux3 mux_904 (.in({n2593, n2582, n2134}), .out(n2154), .config_in(config_chain[6355:6354])); 
mux3 mux_905 (.in({n2707, n2672, n2175}), .out(n2155), .config_in(config_chain[6357:6356])); 
mux3 mux_906 (.in({n2595, n2580, n2136}), .out(n2156), .config_in(config_chain[6359:6358])); 
mux3 mux_907 (.in({n2705, n2674, n2177}), .out(n2157), .config_in(config_chain[6361:6360])); 
mux3 mux_908 (.in({n2597, n2578, n2138}), .out(n2158), .config_in(config_chain[6363:6362])); 
mux3 mux_909 (.in({n2703, n2676, n2179}), .out(n2159), .config_in(config_chain[6365:6364])); 
mux3 mux_910 (.in({n2599, n2576, n2140}), .out(n2160), .config_in(config_chain[6367:6366])); 
mux3 mux_911 (.in({n2701, n2678, n2181}), .out(n2161), .config_in(config_chain[6369:6368])); 
mux3 mux_912 (.in({n2601, n2574, n2142}), .out(n2162), .config_in(config_chain[6371:6370])); 
mux3 mux_913 (.in({n2699, n2680, n2183}), .out(n2163), .config_in(config_chain[6373:6372])); 
mux3 mux_914 (.in({n2603, n2572, n2144}), .out(n2164), .config_in(config_chain[6375:6374])); 
mux3 mux_915 (.in({n2697, n2682, n2185}), .out(n2165), .config_in(config_chain[6377:6376])); 
mux3 mux_916 (.in({n2605, n2570, n2146}), .out(n2166), .config_in(config_chain[6379:6378])); 
mux3 mux_917 (.in({n2695, n2684, n2187}), .out(n2167), .config_in(config_chain[6381:6380])); 
mux3 mux_918 (.in({n2607, n2588, n2148}), .out(n2168), .config_in(config_chain[6383:6382])); 
mux3 mux_919 (.in({n2693, n2686, n2189}), .out(n2169), .config_in(config_chain[6385:6384])); 
mux4 mux_920 (.in({n2709, n2686, n2150, n1143}), .out(n2170), .config_in(config_chain[6387:6386])); 
mux4 mux_921 (.in({n2791, n2788, n2191, n1143}), .out(n2171), .config_in(config_chain[6389:6388])); 
mux4 mux_922 (.in({n2691, n2684, n2152, n1143}), .out(n2172), .config_in(config_chain[6391:6390])); 
mux4 mux_923 (.in({n2809, n2770, n2193, n1143}), .out(n2173), .config_in(config_chain[6393:6392])); 
mux3 mux_924 (.in({n2693, n2682, n2154}), .out(n2174), .config_in(config_chain[6395:6394])); 
mux3 mux_925 (.in({n2807, n2772, n2195}), .out(n2175), .config_in(config_chain[6397:6396])); 
mux3 mux_926 (.in({n2695, n2680, n2156}), .out(n2176), .config_in(config_chain[6399:6398])); 
mux3 mux_927 (.in({n2805, n2774, n2197}), .out(n2177), .config_in(config_chain[6401:6400])); 
mux3 mux_928 (.in({n2697, n2678, n2158}), .out(n2178), .config_in(config_chain[6403:6402])); 
mux3 mux_929 (.in({n2803, n2776, n2199}), .out(n2179), .config_in(config_chain[6405:6404])); 
mux3 mux_930 (.in({n2699, n2676, n2160}), .out(n2180), .config_in(config_chain[6407:6406])); 
mux3 mux_931 (.in({n2801, n2778, n2201}), .out(n2181), .config_in(config_chain[6409:6408])); 
mux3 mux_932 (.in({n2701, n2674, n2162}), .out(n2182), .config_in(config_chain[6411:6410])); 
mux3 mux_933 (.in({n2799, n2780, n2203}), .out(n2183), .config_in(config_chain[6413:6412])); 
mux3 mux_934 (.in({n2703, n2672, n2164}), .out(n2184), .config_in(config_chain[6415:6414])); 
mux3 mux_935 (.in({n2797, n2782, n2205}), .out(n2185), .config_in(config_chain[6417:6416])); 
mux3 mux_936 (.in({n2705, n2670, n2166}), .out(n2186), .config_in(config_chain[6419:6418])); 
mux3 mux_937 (.in({n2795, n2784, n2207}), .out(n2187), .config_in(config_chain[6421:6420])); 
mux3 mux_938 (.in({n2707, n2688, n2168}), .out(n2188), .config_in(config_chain[6423:6422])); 
mux3 mux_939 (.in({n2793, n2786, n2209}), .out(n2189), .config_in(config_chain[6425:6424])); 
mux4 mux_940 (.in({n2809, n2786, n2170, n1389}), .out(n2190), .config_in(config_chain[6427:6426])); 
mux3 mux_941 (.in({n2891, n2870, n1389}), .out(n2191), .config_in(config_chain[6429:6428])); 
mux4 mux_942 (.in({n2791, n2784, n2172, n1389}), .out(n2192), .config_in(config_chain[6431:6430])); 
mux3 mux_943 (.in({n2899, n2878, n1389}), .out(n2193), .config_in(config_chain[6433:6432])); 
mux3 mux_944 (.in({n2793, n2782, n2174}), .out(n2194), .config_in(config_chain[6435:6434])); 
mux2 mux_945 (.in({n2901, n2880}), .out(n2195), .config_in(config_chain[6436:6436])); 
mux3 mux_946 (.in({n2795, n2780, n2176}), .out(n2196), .config_in(config_chain[6438:6437])); 
mux2 mux_947 (.in({n2893, n2872}), .out(n2197), .config_in(config_chain[6439:6439])); 
mux3 mux_948 (.in({n2797, n2778, n2178}), .out(n2198), .config_in(config_chain[6441:6440])); 
mux2 mux_949 (.in({n2903, n2882}), .out(n2199), .config_in(config_chain[6442:6442])); 
mux3 mux_950 (.in({n2799, n2776, n2180}), .out(n2200), .config_in(config_chain[6444:6443])); 
mux2 mux_951 (.in({n2905, n2884}), .out(n2201), .config_in(config_chain[6445:6445])); 
mux3 mux_952 (.in({n2801, n2774, n2182}), .out(n2202), .config_in(config_chain[6447:6446])); 
mux2 mux_953 (.in({n2895, n2874}), .out(n2203), .config_in(config_chain[6448:6448])); 
mux3 mux_954 (.in({n2803, n2772, n2184}), .out(n2204), .config_in(config_chain[6450:6449])); 
mux2 mux_955 (.in({n2907, n2886}), .out(n2205), .config_in(config_chain[6451:6451])); 
mux3 mux_956 (.in({n2805, n2770, n2186}), .out(n2206), .config_in(config_chain[6453:6452])); 
mux2 mux_957 (.in({n2909, n2888}), .out(n2207), .config_in(config_chain[6454:6454])); 
mux3 mux_958 (.in({n2807, n2788, n2188}), .out(n2208), .config_in(config_chain[6456:6455])); 
mux2 mux_959 (.in({n2897, n2876}), .out(n2209), .config_in(config_chain[6457:6457])); 
mux3 mux_960 (.in({n2406, n475, n435}), .out(n2210), .config_in(config_chain[6459:6458])); 
mux4 mux_961 (.in({n2490, n2231, n475, n435}), .out(n2211), .config_in(config_chain[6461:6460])); 
mux3 mux_962 (.in({n2404, n475, n435}), .out(n2212), .config_in(config_chain[6463:6462])); 
mux4 mux_963 (.in({n2492, n2233, n475, n435}), .out(n2213), .config_in(config_chain[6465:6464])); 
mux3 mux_964 (.in({n2402, n478, n463}), .out(n2214), .config_in(config_chain[6467:6466])); 
mux4 mux_965 (.in({n2494, n2235, n478, n463}), .out(n2215), .config_in(config_chain[6469:6468])); 
mux3 mux_966 (.in({n2400, n478, n463}), .out(n2216), .config_in(config_chain[6471:6470])); 
mux4 mux_967 (.in({n2496, n2237, n478, n463}), .out(n2217), .config_in(config_chain[6473:6472])); 
mux3 mux_968 (.in({n2398, n481, n466}), .out(n2218), .config_in(config_chain[6475:6474])); 
mux4 mux_969 (.in({n2498, n2239, n481, n466}), .out(n2219), .config_in(config_chain[6477:6476])); 
mux3 mux_970 (.in({n2396, n481, n466}), .out(n2220), .config_in(config_chain[6479:6478])); 
mux4 mux_971 (.in({n2500, n2241, n481, n466}), .out(n2221), .config_in(config_chain[6481:6480])); 
mux3 mux_972 (.in({n2394, n484, n469}), .out(n2222), .config_in(config_chain[6483:6482])); 
mux4 mux_973 (.in({n2502, n2243, n484, n469}), .out(n2223), .config_in(config_chain[6485:6484])); 
mux3 mux_974 (.in({n2392, n484, n469}), .out(n2224), .config_in(config_chain[6487:6486])); 
mux4 mux_975 (.in({n2504, n2245, n484, n469}), .out(n2225), .config_in(config_chain[6489:6488])); 
mux2 mux_976 (.in({n2390, n472}), .out(n2226), .config_in(config_chain[6490:6490])); 
mux3 mux_977 (.in({n2506, n2247, n472}), .out(n2227), .config_in(config_chain[6492:6491])); 
mux2 mux_978 (.in({n2408, n472}), .out(n2228), .config_in(config_chain[6493:6493])); 
mux3 mux_979 (.in({n2508, n2249, n472}), .out(n2229), .config_in(config_chain[6495:6494])); 
mux4 mux_980 (.in({n2490, n2210, n721, n681}), .out(n2230), .config_in(config_chain[6497:6496])); 
mux4 mux_981 (.in({n2590, n2251, n721, n681}), .out(n2231), .config_in(config_chain[6499:6498])); 
mux4 mux_982 (.in({n2492, n2212, n721, n681}), .out(n2232), .config_in(config_chain[6501:6500])); 
mux4 mux_983 (.in({n2592, n2253, n721, n681}), .out(n2233), .config_in(config_chain[6503:6502])); 
mux4 mux_984 (.in({n2494, n2214, n724, n709}), .out(n2234), .config_in(config_chain[6505:6504])); 
mux4 mux_985 (.in({n2594, n2255, n724, n709}), .out(n2235), .config_in(config_chain[6507:6506])); 
mux4 mux_986 (.in({n2496, n2216, n724, n709}), .out(n2236), .config_in(config_chain[6509:6508])); 
mux4 mux_987 (.in({n2596, n2257, n724, n709}), .out(n2237), .config_in(config_chain[6511:6510])); 
mux4 mux_988 (.in({n2498, n2218, n727, n712}), .out(n2238), .config_in(config_chain[6513:6512])); 
mux4 mux_989 (.in({n2598, n2259, n727, n712}), .out(n2239), .config_in(config_chain[6515:6514])); 
mux4 mux_990 (.in({n2500, n2220, n727, n712}), .out(n2240), .config_in(config_chain[6517:6516])); 
mux4 mux_991 (.in({n2600, n2261, n727, n712}), .out(n2241), .config_in(config_chain[6519:6518])); 
mux4 mux_992 (.in({n2502, n2222, n730, n715}), .out(n2242), .config_in(config_chain[6521:6520])); 
mux4 mux_993 (.in({n2602, n2263, n730, n715}), .out(n2243), .config_in(config_chain[6523:6522])); 
mux4 mux_994 (.in({n2504, n2224, n730, n715}), .out(n2244), .config_in(config_chain[6525:6524])); 
mux4 mux_995 (.in({n2604, n2265, n730, n715}), .out(n2245), .config_in(config_chain[6527:6526])); 
mux3 mux_996 (.in({n2506, n2226, n718}), .out(n2246), .config_in(config_chain[6529:6528])); 
mux3 mux_997 (.in({n2606, n2267, n718}), .out(n2247), .config_in(config_chain[6531:6530])); 
mux3 mux_998 (.in({n2508, n2228, n718}), .out(n2248), .config_in(config_chain[6533:6532])); 
mux3 mux_999 (.in({n2608, n2269, n718}), .out(n2249), .config_in(config_chain[6535:6534])); 
mux4 mux_1000 (.in({n2590, n2230, n967, n927}), .out(n2250), .config_in(config_chain[6537:6536])); 
mux4 mux_1001 (.in({n2690, n2271, n967, n927}), .out(n2251), .config_in(config_chain[6539:6538])); 
mux4 mux_1002 (.in({n2592, n2232, n967, n927}), .out(n2252), .config_in(config_chain[6541:6540])); 
mux4 mux_1003 (.in({n2692, n2273, n967, n927}), .out(n2253), .config_in(config_chain[6543:6542])); 
mux4 mux_1004 (.in({n2594, n2234, n970, n955}), .out(n2254), .config_in(config_chain[6545:6544])); 
mux4 mux_1005 (.in({n2694, n2275, n970, n955}), .out(n2255), .config_in(config_chain[6547:6546])); 
mux4 mux_1006 (.in({n2596, n2236, n970, n955}), .out(n2256), .config_in(config_chain[6549:6548])); 
mux4 mux_1007 (.in({n2696, n2277, n970, n955}), .out(n2257), .config_in(config_chain[6551:6550])); 
mux4 mux_1008 (.in({n2598, n2238, n973, n958}), .out(n2258), .config_in(config_chain[6553:6552])); 
mux4 mux_1009 (.in({n2698, n2279, n973, n958}), .out(n2259), .config_in(config_chain[6555:6554])); 
mux4 mux_1010 (.in({n2600, n2240, n973, n958}), .out(n2260), .config_in(config_chain[6557:6556])); 
mux4 mux_1011 (.in({n2700, n2281, n973, n958}), .out(n2261), .config_in(config_chain[6559:6558])); 
mux4 mux_1012 (.in({n2602, n2242, n976, n961}), .out(n2262), .config_in(config_chain[6561:6560])); 
mux4 mux_1013 (.in({n2702, n2283, n976, n961}), .out(n2263), .config_in(config_chain[6563:6562])); 
mux4 mux_1014 (.in({n2604, n2244, n976, n961}), .out(n2264), .config_in(config_chain[6565:6564])); 
mux4 mux_1015 (.in({n2704, n2285, n976, n961}), .out(n2265), .config_in(config_chain[6567:6566])); 
mux3 mux_1016 (.in({n2606, n2246, n964}), .out(n2266), .config_in(config_chain[6569:6568])); 
mux3 mux_1017 (.in({n2706, n2287, n964}), .out(n2267), .config_in(config_chain[6571:6570])); 
mux3 mux_1018 (.in({n2608, n2248, n964}), .out(n2268), .config_in(config_chain[6573:6572])); 
mux3 mux_1019 (.in({n2708, n2289, n964}), .out(n2269), .config_in(config_chain[6575:6574])); 
mux4 mux_1020 (.in({n2690, n2250, n1213, n1173}), .out(n2270), .config_in(config_chain[6577:6576])); 
mux4 mux_1021 (.in({n2790, n2291, n1213, n1173}), .out(n2271), .config_in(config_chain[6579:6578])); 
mux4 mux_1022 (.in({n2692, n2252, n1213, n1173}), .out(n2272), .config_in(config_chain[6581:6580])); 
mux4 mux_1023 (.in({n2792, n2293, n1213, n1173}), .out(n2273), .config_in(config_chain[6583:6582])); 
mux4 mux_1024 (.in({n2694, n2254, n1216, n1201}), .out(n2274), .config_in(config_chain[6585:6584])); 
mux4 mux_1025 (.in({n2794, n2295, n1216, n1201}), .out(n2275), .config_in(config_chain[6587:6586])); 
mux4 mux_1026 (.in({n2696, n2256, n1216, n1201}), .out(n2276), .config_in(config_chain[6589:6588])); 
mux4 mux_1027 (.in({n2796, n2297, n1216, n1201}), .out(n2277), .config_in(config_chain[6591:6590])); 
mux4 mux_1028 (.in({n2698, n2258, n1219, n1204}), .out(n2278), .config_in(config_chain[6593:6592])); 
mux4 mux_1029 (.in({n2798, n2299, n1219, n1204}), .out(n2279), .config_in(config_chain[6595:6594])); 
mux4 mux_1030 (.in({n2700, n2260, n1219, n1204}), .out(n2280), .config_in(config_chain[6597:6596])); 
mux4 mux_1031 (.in({n2800, n2301, n1219, n1204}), .out(n2281), .config_in(config_chain[6599:6598])); 
mux4 mux_1032 (.in({n2702, n2262, n1222, n1207}), .out(n2282), .config_in(config_chain[6601:6600])); 
mux4 mux_1033 (.in({n2802, n2303, n1222, n1207}), .out(n2283), .config_in(config_chain[6603:6602])); 
mux4 mux_1034 (.in({n2704, n2264, n1222, n1207}), .out(n2284), .config_in(config_chain[6605:6604])); 
mux4 mux_1035 (.in({n2804, n2305, n1222, n1207}), .out(n2285), .config_in(config_chain[6607:6606])); 
mux3 mux_1036 (.in({n2706, n2266, n1210}), .out(n2286), .config_in(config_chain[6609:6608])); 
mux3 mux_1037 (.in({n2806, n2307, n1210}), .out(n2287), .config_in(config_chain[6611:6610])); 
mux3 mux_1038 (.in({n2708, n2268, n1210}), .out(n2288), .config_in(config_chain[6613:6612])); 
mux3 mux_1039 (.in({n2808, n2309, n1210}), .out(n2289), .config_in(config_chain[6615:6614])); 
mux4 mux_1040 (.in({n2790, n2270, n1459, n1419}), .out(n2290), .config_in(config_chain[6617:6616])); 
mux3 mux_1041 (.in({n2908, n1459, n1419}), .out(n2291), .config_in(config_chain[6619:6618])); 
mux4 mux_1042 (.in({n2792, n2272, n1459, n1419}), .out(n2292), .config_in(config_chain[6621:6620])); 
mux3 mux_1043 (.in({n2890, n1459, n1419}), .out(n2293), .config_in(config_chain[6623:6622])); 
mux4 mux_1044 (.in({n2794, n2274, n1462, n1447}), .out(n2294), .config_in(config_chain[6625:6624])); 
mux3 mux_1045 (.in({n2892, n1462, n1447}), .out(n2295), .config_in(config_chain[6627:6626])); 
mux4 mux_1046 (.in({n2796, n2276, n1462, n1447}), .out(n2296), .config_in(config_chain[6629:6628])); 
mux3 mux_1047 (.in({n2894, n1462, n1447}), .out(n2297), .config_in(config_chain[6631:6630])); 
mux4 mux_1048 (.in({n2798, n2278, n1465, n1450}), .out(n2298), .config_in(config_chain[6633:6632])); 
mux3 mux_1049 (.in({n2896, n1465, n1450}), .out(n2299), .config_in(config_chain[6635:6634])); 
mux4 mux_1050 (.in({n2800, n2280, n1465, n1450}), .out(n2300), .config_in(config_chain[6637:6636])); 
mux3 mux_1051 (.in({n2898, n1465, n1450}), .out(n2301), .config_in(config_chain[6639:6638])); 
mux4 mux_1052 (.in({n2802, n2282, n1468, n1453}), .out(n2302), .config_in(config_chain[6641:6640])); 
mux3 mux_1053 (.in({n2900, n1468, n1453}), .out(n2303), .config_in(config_chain[6643:6642])); 
mux4 mux_1054 (.in({n2804, n2284, n1468, n1453}), .out(n2304), .config_in(config_chain[6645:6644])); 
mux3 mux_1055 (.in({n2902, n1468, n1453}), .out(n2305), .config_in(config_chain[6647:6646])); 
mux3 mux_1056 (.in({n2806, n2286, n1456}), .out(n2306), .config_in(config_chain[6649:6648])); 
mux2 mux_1057 (.in({n2904, n1456}), .out(n2307), .config_in(config_chain[6650:6650])); 
mux3 mux_1058 (.in({n2808, n2288, n1456}), .out(n2308), .config_in(config_chain[6652:6651])); 
mux2 mux_1059 (.in({n2906, n1456}), .out(n2309), .config_in(config_chain[6653:6653])); 
mux3 mux_1060 (.in({n1713, n40, n25}), .out(n2310), .config_in(config_chain[6655:6654])); 
mux4 mux_1061 (.in({n2331, n1811, n40, n25}), .out(n2311), .config_in(config_chain[6657:6656])); 
mux3 mux_1062 (.in({n1715, n40, n25}), .out(n2312), .config_in(config_chain[6659:6658])); 
mux4 mux_1063 (.in({n2333, n1813, n40, n25}), .out(n2313), .config_in(config_chain[6661:6660])); 
mux3 mux_1064 (.in({n1717, n43, n28}), .out(n2314), .config_in(config_chain[6663:6662])); 
mux4 mux_1065 (.in({n2335, n1815, n43, n28}), .out(n2315), .config_in(config_chain[6665:6664])); 
mux3 mux_1066 (.in({n1719, n43, n28}), .out(n2316), .config_in(config_chain[6667:6666])); 
mux4 mux_1067 (.in({n2337, n1817, n43, n28}), .out(n2317), .config_in(config_chain[6669:6668])); 
mux3 mux_1068 (.in({n1721, n46, n31}), .out(n2318), .config_in(config_chain[6671:6670])); 
mux4 mux_1069 (.in({n2339, n1819, n46, n31}), .out(n2319), .config_in(config_chain[6673:6672])); 
mux3 mux_1070 (.in({n1723, n46, n31}), .out(n2320), .config_in(config_chain[6675:6674])); 
mux4 mux_1071 (.in({n2341, n1821, n46, n31}), .out(n2321), .config_in(config_chain[6677:6676])); 
mux2 mux_1072 (.in({n1725, n34}), .out(n2322), .config_in(config_chain[6678:6678])); 
mux3 mux_1073 (.in({n2343, n1823, n34}), .out(n2323), .config_in(config_chain[6680:6679])); 
mux2 mux_1074 (.in({n1727, n34}), .out(n2324), .config_in(config_chain[6681:6681])); 
mux3 mux_1075 (.in({n2345, n1825, n34}), .out(n2325), .config_in(config_chain[6683:6682])); 
mux2 mux_1076 (.in({n1729, n37}), .out(n2326), .config_in(config_chain[6684:6684])); 
mux3 mux_1077 (.in({n2347, n1827, n37}), .out(n2327), .config_in(config_chain[6686:6685])); 
mux2 mux_1078 (.in({n1711, n37}), .out(n2328), .config_in(config_chain[6687:6687])); 
mux3 mux_1079 (.in({n2349, n1829, n37}), .out(n2329), .config_in(config_chain[6689:6688])); 
mux4 mux_1080 (.in({n2310, n1811, n88, n73}), .out(n2330), .config_in(config_chain[6691:6690])); 
mux4 mux_1081 (.in({n2351, n1911, n88, n73}), .out(n2331), .config_in(config_chain[6693:6692])); 
mux4 mux_1082 (.in({n2312, n1813, n88, n73}), .out(n2332), .config_in(config_chain[6695:6694])); 
mux4 mux_1083 (.in({n2353, n1913, n88, n73}), .out(n2333), .config_in(config_chain[6697:6696])); 
mux4 mux_1084 (.in({n2314, n1815, n91, n76}), .out(n2334), .config_in(config_chain[6699:6698])); 
mux4 mux_1085 (.in({n2355, n1915, n91, n76}), .out(n2335), .config_in(config_chain[6701:6700])); 
mux4 mux_1086 (.in({n2316, n1817, n91, n76}), .out(n2336), .config_in(config_chain[6703:6702])); 
mux4 mux_1087 (.in({n2357, n1917, n91, n76}), .out(n2337), .config_in(config_chain[6705:6704])); 
mux4 mux_1088 (.in({n2318, n1819, n94, n79}), .out(n2338), .config_in(config_chain[6707:6706])); 
mux4 mux_1089 (.in({n2359, n1919, n94, n79}), .out(n2339), .config_in(config_chain[6709:6708])); 
mux4 mux_1090 (.in({n2320, n1821, n94, n79}), .out(n2340), .config_in(config_chain[6711:6710])); 
mux4 mux_1091 (.in({n2361, n1921, n94, n79}), .out(n2341), .config_in(config_chain[6713:6712])); 
mux3 mux_1092 (.in({n2322, n1823, n82}), .out(n2342), .config_in(config_chain[6715:6714])); 
mux3 mux_1093 (.in({n2363, n1923, n82}), .out(n2343), .config_in(config_chain[6717:6716])); 
mux3 mux_1094 (.in({n2324, n1825, n82}), .out(n2344), .config_in(config_chain[6719:6718])); 
mux3 mux_1095 (.in({n2365, n1925, n82}), .out(n2345), .config_in(config_chain[6721:6720])); 
mux3 mux_1096 (.in({n2326, n1827, n85}), .out(n2346), .config_in(config_chain[6723:6722])); 
mux3 mux_1097 (.in({n2367, n1927, n85}), .out(n2347), .config_in(config_chain[6725:6724])); 
mux3 mux_1098 (.in({n2328, n1829, n85}), .out(n2348), .config_in(config_chain[6727:6726])); 
mux3 mux_1099 (.in({n2369, n1929, n85}), .out(n2349), .config_in(config_chain[6729:6728])); 
mux4 mux_1100 (.in({n2330, n1911, n136, n121}), .out(n2350), .config_in(config_chain[6731:6730])); 
mux4 mux_1101 (.in({n2371, n2011, n136, n121}), .out(n2351), .config_in(config_chain[6733:6732])); 
mux4 mux_1102 (.in({n2332, n1913, n136, n121}), .out(n2352), .config_in(config_chain[6735:6734])); 
mux4 mux_1103 (.in({n2373, n2013, n136, n121}), .out(n2353), .config_in(config_chain[6737:6736])); 
mux4 mux_1104 (.in({n2334, n1915, n139, n124}), .out(n2354), .config_in(config_chain[6739:6738])); 
mux4 mux_1105 (.in({n2375, n2015, n139, n124}), .out(n2355), .config_in(config_chain[6741:6740])); 
mux4 mux_1106 (.in({n2336, n1917, n139, n124}), .out(n2356), .config_in(config_chain[6743:6742])); 
mux4 mux_1107 (.in({n2377, n2017, n139, n124}), .out(n2357), .config_in(config_chain[6745:6744])); 
mux4 mux_1108 (.in({n2338, n1919, n142, n127}), .out(n2358), .config_in(config_chain[6747:6746])); 
mux4 mux_1109 (.in({n2379, n2019, n142, n127}), .out(n2359), .config_in(config_chain[6749:6748])); 
mux4 mux_1110 (.in({n2340, n1921, n142, n127}), .out(n2360), .config_in(config_chain[6751:6750])); 
mux4 mux_1111 (.in({n2381, n2021, n142, n127}), .out(n2361), .config_in(config_chain[6753:6752])); 
mux3 mux_1112 (.in({n2342, n1923, n130}), .out(n2362), .config_in(config_chain[6755:6754])); 
mux3 mux_1113 (.in({n2383, n2023, n130}), .out(n2363), .config_in(config_chain[6757:6756])); 
mux3 mux_1114 (.in({n2344, n1925, n130}), .out(n2364), .config_in(config_chain[6759:6758])); 
mux3 mux_1115 (.in({n2385, n2025, n130}), .out(n2365), .config_in(config_chain[6761:6760])); 
mux3 mux_1116 (.in({n2346, n1927, n133}), .out(n2366), .config_in(config_chain[6763:6762])); 
mux3 mux_1117 (.in({n2387, n2027, n133}), .out(n2367), .config_in(config_chain[6765:6764])); 
mux3 mux_1118 (.in({n2348, n1929, n133}), .out(n2368), .config_in(config_chain[6767:6766])); 
mux3 mux_1119 (.in({n2389, n2029, n133}), .out(n2369), .config_in(config_chain[6769:6768])); 
mux4 mux_1120 (.in({n2350, n2011, n184, n169}), .out(n2370), .config_in(config_chain[6771:6770])); 
mux4 mux_1121 (.in({n2391, n2111, n184, n169}), .out(n2371), .config_in(config_chain[6773:6772])); 
mux4 mux_1122 (.in({n2352, n2013, n184, n169}), .out(n2372), .config_in(config_chain[6775:6774])); 
mux4 mux_1123 (.in({n2393, n2113, n184, n169}), .out(n2373), .config_in(config_chain[6777:6776])); 
mux4 mux_1124 (.in({n2354, n2015, n187, n172}), .out(n2374), .config_in(config_chain[6779:6778])); 
mux4 mux_1125 (.in({n2395, n2115, n187, n172}), .out(n2375), .config_in(config_chain[6781:6780])); 
mux4 mux_1126 (.in({n2356, n2017, n187, n172}), .out(n2376), .config_in(config_chain[6783:6782])); 
mux4 mux_1127 (.in({n2397, n2117, n187, n172}), .out(n2377), .config_in(config_chain[6785:6784])); 
mux4 mux_1128 (.in({n2358, n2019, n190, n175}), .out(n2378), .config_in(config_chain[6787:6786])); 
mux4 mux_1129 (.in({n2399, n2119, n190, n175}), .out(n2379), .config_in(config_chain[6789:6788])); 
mux4 mux_1130 (.in({n2360, n2021, n190, n175}), .out(n2380), .config_in(config_chain[6791:6790])); 
mux4 mux_1131 (.in({n2401, n2121, n190, n175}), .out(n2381), .config_in(config_chain[6793:6792])); 
mux3 mux_1132 (.in({n2362, n2023, n178}), .out(n2382), .config_in(config_chain[6795:6794])); 
mux3 mux_1133 (.in({n2403, n2123, n178}), .out(n2383), .config_in(config_chain[6797:6796])); 
mux3 mux_1134 (.in({n2364, n2025, n178}), .out(n2384), .config_in(config_chain[6799:6798])); 
mux3 mux_1135 (.in({n2405, n2125, n178}), .out(n2385), .config_in(config_chain[6801:6800])); 
mux3 mux_1136 (.in({n2366, n2027, n181}), .out(n2386), .config_in(config_chain[6803:6802])); 
mux3 mux_1137 (.in({n2407, n2127, n181}), .out(n2387), .config_in(config_chain[6805:6804])); 
mux3 mux_1138 (.in({n2368, n2029, n181}), .out(n2388), .config_in(config_chain[6807:6806])); 
mux3 mux_1139 (.in({n2409, n2129, n181}), .out(n2389), .config_in(config_chain[6809:6808])); 
mux4 mux_1140 (.in({n2370, n2111, n232, n217}), .out(n2390), .config_in(config_chain[6811:6810])); 
mux3 mux_1141 (.in({n2227, n232, n217}), .out(n2391), .config_in(config_chain[6813:6812])); 
mux4 mux_1142 (.in({n2372, n2113, n232, n217}), .out(n2392), .config_in(config_chain[6815:6814])); 
mux3 mux_1143 (.in({n2225, n232, n217}), .out(n2393), .config_in(config_chain[6817:6816])); 
mux4 mux_1144 (.in({n2374, n2115, n235, n220}), .out(n2394), .config_in(config_chain[6819:6818])); 
mux3 mux_1145 (.in({n2223, n235, n220}), .out(n2395), .config_in(config_chain[6821:6820])); 
mux4 mux_1146 (.in({n2376, n2117, n235, n220}), .out(n2396), .config_in(config_chain[6823:6822])); 
mux3 mux_1147 (.in({n2221, n235, n220}), .out(n2397), .config_in(config_chain[6825:6824])); 
mux4 mux_1148 (.in({n2378, n2119, n238, n223}), .out(n2398), .config_in(config_chain[6827:6826])); 
mux3 mux_1149 (.in({n2219, n238, n223}), .out(n2399), .config_in(config_chain[6829:6828])); 
mux4 mux_1150 (.in({n2380, n2121, n238, n223}), .out(n2400), .config_in(config_chain[6831:6830])); 
mux3 mux_1151 (.in({n2217, n238, n223}), .out(n2401), .config_in(config_chain[6833:6832])); 
mux3 mux_1152 (.in({n2382, n2123, n226}), .out(n2402), .config_in(config_chain[6835:6834])); 
mux2 mux_1153 (.in({n2215, n226}), .out(n2403), .config_in(config_chain[6836:6836])); 
mux3 mux_1154 (.in({n2384, n2125, n226}), .out(n2404), .config_in(config_chain[6838:6837])); 
mux2 mux_1155 (.in({n2213, n226}), .out(n2405), .config_in(config_chain[6839:6839])); 
mux3 mux_1156 (.in({n2386, n2127, n229}), .out(n2406), .config_in(config_chain[6841:6840])); 
mux2 mux_1157 (.in({n2211, n229}), .out(n2407), .config_in(config_chain[6842:6842])); 
mux3 mux_1158 (.in({n2388, n2129, n229}), .out(n2408), .config_in(config_chain[6844:6843])); 
mux2 mux_1159 (.in({n2229, n229}), .out(n2409), .config_in(config_chain[6845:6845])); 
mux3 mux_1160 (.in({n1737, n1716, n316}), .out(n2410), .config_in(config_chain[6847:6846])); 
mux4 mux_1161 (.in({n2431, n1847, n1812, n316}), .out(n2411), .config_in(config_chain[6849:6848])); 
mux3 mux_1162 (.in({n1739, n1718, n316}), .out(n2412), .config_in(config_chain[6851:6850])); 
mux4 mux_1163 (.in({n2433, n1845, n1814, n316}), .out(n2413), .config_in(config_chain[6853:6852])); 
mux2 mux_1164 (.in({n1731, n1710}), .out(n2414), .config_in(config_chain[6854:6854])); 
mux3 mux_1165 (.in({n2435, n1843, n1816}), .out(n2415), .config_in(config_chain[6856:6855])); 
mux2 mux_1166 (.in({n1741, n1720}), .out(n2416), .config_in(config_chain[6857:6857])); 
mux3 mux_1167 (.in({n2437, n1841, n1818}), .out(n2417), .config_in(config_chain[6859:6858])); 
mux2 mux_1168 (.in({n1743, n1722}), .out(n2418), .config_in(config_chain[6860:6860])); 
mux3 mux_1169 (.in({n2439, n1839, n1820}), .out(n2419), .config_in(config_chain[6862:6861])); 
mux2 mux_1170 (.in({n1733, n1712}), .out(n2420), .config_in(config_chain[6863:6863])); 
mux3 mux_1171 (.in({n2441, n1837, n1822}), .out(n2421), .config_in(config_chain[6865:6864])); 
mux2 mux_1172 (.in({n1745, n1724}), .out(n2422), .config_in(config_chain[6866:6866])); 
mux3 mux_1173 (.in({n2443, n1835, n1824}), .out(n2423), .config_in(config_chain[6868:6867])); 
mux2 mux_1174 (.in({n1747, n1726}), .out(n2424), .config_in(config_chain[6869:6869])); 
mux3 mux_1175 (.in({n2445, n1833, n1826}), .out(n2425), .config_in(config_chain[6871:6870])); 
mux2 mux_1176 (.in({n1735, n1714}), .out(n2426), .config_in(config_chain[6872:6872])); 
mux3 mux_1177 (.in({n2447, n1831, n1828}), .out(n2427), .config_in(config_chain[6874:6873])); 
mux2 mux_1178 (.in({n1749, n1728}), .out(n2428), .config_in(config_chain[6875:6875])); 
mux3 mux_1179 (.in({n2449, n1849, n1810}), .out(n2429), .config_in(config_chain[6877:6876])); 
mux4 mux_1180 (.in({n2410, n1833, n1810, n346}), .out(n2430), .config_in(config_chain[6879:6878])); 
mux4 mux_1181 (.in({n2451, n1947, n1912, n346}), .out(n2431), .config_in(config_chain[6881:6880])); 
mux4 mux_1182 (.in({n2412, n1835, n1828, n346}), .out(n2432), .config_in(config_chain[6883:6882])); 
mux4 mux_1183 (.in({n2453, n1945, n1914, n346}), .out(n2433), .config_in(config_chain[6885:6884])); 
mux3 mux_1184 (.in({n2414, n1837, n1826}), .out(n2434), .config_in(config_chain[6887:6886])); 
mux3 mux_1185 (.in({n2455, n1943, n1916}), .out(n2435), .config_in(config_chain[6889:6888])); 
mux3 mux_1186 (.in({n2416, n1839, n1824}), .out(n2436), .config_in(config_chain[6891:6890])); 
mux3 mux_1187 (.in({n2457, n1941, n1918}), .out(n2437), .config_in(config_chain[6893:6892])); 
mux3 mux_1188 (.in({n2418, n1841, n1822}), .out(n2438), .config_in(config_chain[6895:6894])); 
mux3 mux_1189 (.in({n2459, n1939, n1920}), .out(n2439), .config_in(config_chain[6897:6896])); 
mux3 mux_1190 (.in({n2420, n1843, n1820}), .out(n2440), .config_in(config_chain[6899:6898])); 
mux3 mux_1191 (.in({n2461, n1937, n1922}), .out(n2441), .config_in(config_chain[6901:6900])); 
mux3 mux_1192 (.in({n2422, n1845, n1818}), .out(n2442), .config_in(config_chain[6903:6902])); 
mux3 mux_1193 (.in({n2463, n1935, n1924}), .out(n2443), .config_in(config_chain[6905:6904])); 
mux3 mux_1194 (.in({n2424, n1847, n1816}), .out(n2444), .config_in(config_chain[6907:6906])); 
mux3 mux_1195 (.in({n2465, n1933, n1926}), .out(n2445), .config_in(config_chain[6909:6908])); 
mux3 mux_1196 (.in({n2426, n1849, n1814}), .out(n2446), .config_in(config_chain[6911:6910])); 
mux3 mux_1197 (.in({n2467, n1931, n1928}), .out(n2447), .config_in(config_chain[6913:6912])); 
mux3 mux_1198 (.in({n2428, n1831, n1812}), .out(n2448), .config_in(config_chain[6915:6914])); 
mux3 mux_1199 (.in({n2469, n1949, n1910}), .out(n2449), .config_in(config_chain[6917:6916])); 
mux4 mux_1200 (.in({n2430, n1933, n1910, n376}), .out(n2450), .config_in(config_chain[6919:6918])); 
mux4 mux_1201 (.in({n2471, n2047, n2012, n376}), .out(n2451), .config_in(config_chain[6921:6920])); 
mux4 mux_1202 (.in({n2432, n1935, n1928, n376}), .out(n2452), .config_in(config_chain[6923:6922])); 
mux4 mux_1203 (.in({n2473, n2045, n2014, n376}), .out(n2453), .config_in(config_chain[6925:6924])); 
mux3 mux_1204 (.in({n2434, n1937, n1926}), .out(n2454), .config_in(config_chain[6927:6926])); 
mux3 mux_1205 (.in({n2475, n2043, n2016}), .out(n2455), .config_in(config_chain[6929:6928])); 
mux3 mux_1206 (.in({n2436, n1939, n1924}), .out(n2456), .config_in(config_chain[6931:6930])); 
mux3 mux_1207 (.in({n2477, n2041, n2018}), .out(n2457), .config_in(config_chain[6933:6932])); 
mux3 mux_1208 (.in({n2438, n1941, n1922}), .out(n2458), .config_in(config_chain[6935:6934])); 
mux3 mux_1209 (.in({n2479, n2039, n2020}), .out(n2459), .config_in(config_chain[6937:6936])); 
mux3 mux_1210 (.in({n2440, n1943, n1920}), .out(n2460), .config_in(config_chain[6939:6938])); 
mux3 mux_1211 (.in({n2481, n2037, n2022}), .out(n2461), .config_in(config_chain[6941:6940])); 
mux3 mux_1212 (.in({n2442, n1945, n1918}), .out(n2462), .config_in(config_chain[6943:6942])); 
mux3 mux_1213 (.in({n2483, n2035, n2024}), .out(n2463), .config_in(config_chain[6945:6944])); 
mux3 mux_1214 (.in({n2444, n1947, n1916}), .out(n2464), .config_in(config_chain[6947:6946])); 
mux3 mux_1215 (.in({n2485, n2033, n2026}), .out(n2465), .config_in(config_chain[6949:6948])); 
mux3 mux_1216 (.in({n2446, n1949, n1914}), .out(n2466), .config_in(config_chain[6951:6950])); 
mux3 mux_1217 (.in({n2487, n2031, n2028}), .out(n2467), .config_in(config_chain[6953:6952])); 
mux3 mux_1218 (.in({n2448, n1931, n1912}), .out(n2468), .config_in(config_chain[6955:6954])); 
mux3 mux_1219 (.in({n2489, n2049, n2010}), .out(n2469), .config_in(config_chain[6957:6956])); 
mux4 mux_1220 (.in({n2450, n2033, n2010, n406}), .out(n2470), .config_in(config_chain[6959:6958])); 
mux4 mux_1221 (.in({n2491, n2147, n2112, n406}), .out(n2471), .config_in(config_chain[6961:6960])); 
mux4 mux_1222 (.in({n2452, n2035, n2028, n406}), .out(n2472), .config_in(config_chain[6963:6962])); 
mux4 mux_1223 (.in({n2493, n2145, n2114, n406}), .out(n2473), .config_in(config_chain[6965:6964])); 
mux3 mux_1224 (.in({n2454, n2037, n2026}), .out(n2474), .config_in(config_chain[6967:6966])); 
mux3 mux_1225 (.in({n2495, n2143, n2116}), .out(n2475), .config_in(config_chain[6969:6968])); 
mux3 mux_1226 (.in({n2456, n2039, n2024}), .out(n2476), .config_in(config_chain[6971:6970])); 
mux3 mux_1227 (.in({n2497, n2141, n2118}), .out(n2477), .config_in(config_chain[6973:6972])); 
mux3 mux_1228 (.in({n2458, n2041, n2022}), .out(n2478), .config_in(config_chain[6975:6974])); 
mux3 mux_1229 (.in({n2499, n2139, n2120}), .out(n2479), .config_in(config_chain[6977:6976])); 
mux3 mux_1230 (.in({n2460, n2043, n2020}), .out(n2480), .config_in(config_chain[6979:6978])); 
mux3 mux_1231 (.in({n2501, n2137, n2122}), .out(n2481), .config_in(config_chain[6981:6980])); 
mux3 mux_1232 (.in({n2462, n2045, n2018}), .out(n2482), .config_in(config_chain[6983:6982])); 
mux3 mux_1233 (.in({n2503, n2135, n2124}), .out(n2483), .config_in(config_chain[6985:6984])); 
mux3 mux_1234 (.in({n2464, n2047, n2016}), .out(n2484), .config_in(config_chain[6987:6986])); 
mux3 mux_1235 (.in({n2505, n2133, n2126}), .out(n2485), .config_in(config_chain[6989:6988])); 
mux3 mux_1236 (.in({n2466, n2049, n2014}), .out(n2486), .config_in(config_chain[6991:6990])); 
mux3 mux_1237 (.in({n2507, n2131, n2128}), .out(n2487), .config_in(config_chain[6993:6992])); 
mux3 mux_1238 (.in({n2468, n2031, n2012}), .out(n2488), .config_in(config_chain[6995:6994])); 
mux3 mux_1239 (.in({n2509, n2149, n2110}), .out(n2489), .config_in(config_chain[6997:6996])); 
mux4 mux_1240 (.in({n2470, n2133, n2110, n436}), .out(n2490), .config_in(config_chain[6999:6998])); 
mux3 mux_1241 (.in({n2231, n2210, n436}), .out(n2491), .config_in(config_chain[7001:7000])); 
mux4 mux_1242 (.in({n2472, n2135, n2128, n436}), .out(n2492), .config_in(config_chain[7003:7002])); 
mux3 mux_1243 (.in({n2239, n2218, n436}), .out(n2493), .config_in(config_chain[7005:7004])); 
mux3 mux_1244 (.in({n2474, n2137, n2126}), .out(n2494), .config_in(config_chain[7007:7006])); 
mux2 mux_1245 (.in({n2241, n2220}), .out(n2495), .config_in(config_chain[7008:7008])); 
mux3 mux_1246 (.in({n2476, n2139, n2124}), .out(n2496), .config_in(config_chain[7010:7009])); 
mux2 mux_1247 (.in({n2233, n2212}), .out(n2497), .config_in(config_chain[7011:7011])); 
mux3 mux_1248 (.in({n2478, n2141, n2122}), .out(n2498), .config_in(config_chain[7013:7012])); 
mux2 mux_1249 (.in({n2243, n2222}), .out(n2499), .config_in(config_chain[7014:7014])); 
mux3 mux_1250 (.in({n2480, n2143, n2120}), .out(n2500), .config_in(config_chain[7016:7015])); 
mux2 mux_1251 (.in({n2245, n2224}), .out(n2501), .config_in(config_chain[7017:7017])); 
mux3 mux_1252 (.in({n2482, n2145, n2118}), .out(n2502), .config_in(config_chain[7019:7018])); 
mux2 mux_1253 (.in({n2235, n2214}), .out(n2503), .config_in(config_chain[7020:7020])); 
mux3 mux_1254 (.in({n2484, n2147, n2116}), .out(n2504), .config_in(config_chain[7022:7021])); 
mux2 mux_1255 (.in({n2247, n2226}), .out(n2505), .config_in(config_chain[7023:7023])); 
mux3 mux_1256 (.in({n2486, n2149, n2114}), .out(n2506), .config_in(config_chain[7025:7024])); 
mux2 mux_1257 (.in({n2249, n2228}), .out(n2507), .config_in(config_chain[7026:7026])); 
mux3 mux_1258 (.in({n2488, n2131, n2112}), .out(n2508), .config_in(config_chain[7028:7027])); 
mux2 mux_1259 (.in({n2237, n2216}), .out(n2509), .config_in(config_chain[7029:7029])); 
mux3 mux_1260 (.in({n1757, n1736, n562}), .out(n2510), .config_in(config_chain[7031:7030])); 
mux4 mux_1261 (.in({n2531, n1867, n1832, n562}), .out(n2511), .config_in(config_chain[7033:7032])); 
mux3 mux_1262 (.in({n1759, n1738, n562}), .out(n2512), .config_in(config_chain[7035:7034])); 
mux4 mux_1263 (.in({n2533, n1865, n1834, n562}), .out(n2513), .config_in(config_chain[7037:7036])); 
mux2 mux_1264 (.in({n1751, n1730}), .out(n2514), .config_in(config_chain[7038:7038])); 
mux3 mux_1265 (.in({n2535, n1863, n1836}), .out(n2515), .config_in(config_chain[7040:7039])); 
mux2 mux_1266 (.in({n1761, n1740}), .out(n2516), .config_in(config_chain[7041:7041])); 
mux3 mux_1267 (.in({n2537, n1861, n1838}), .out(n2517), .config_in(config_chain[7043:7042])); 
mux2 mux_1268 (.in({n1763, n1742}), .out(n2518), .config_in(config_chain[7044:7044])); 
mux3 mux_1269 (.in({n2539, n1859, n1840}), .out(n2519), .config_in(config_chain[7046:7045])); 
mux2 mux_1270 (.in({n1753, n1732}), .out(n2520), .config_in(config_chain[7047:7047])); 
mux3 mux_1271 (.in({n2541, n1857, n1842}), .out(n2521), .config_in(config_chain[7049:7048])); 
mux2 mux_1272 (.in({n1765, n1744}), .out(n2522), .config_in(config_chain[7050:7050])); 
mux3 mux_1273 (.in({n2543, n1855, n1844}), .out(n2523), .config_in(config_chain[7052:7051])); 
mux2 mux_1274 (.in({n1767, n1746}), .out(n2524), .config_in(config_chain[7053:7053])); 
mux3 mux_1275 (.in({n2545, n1853, n1846}), .out(n2525), .config_in(config_chain[7055:7054])); 
mux2 mux_1276 (.in({n1755, n1734}), .out(n2526), .config_in(config_chain[7056:7056])); 
mux3 mux_1277 (.in({n2547, n1851, n1848}), .out(n2527), .config_in(config_chain[7058:7057])); 
mux2 mux_1278 (.in({n1769, n1748}), .out(n2528), .config_in(config_chain[7059:7059])); 
mux3 mux_1279 (.in({n2549, n1869, n1830}), .out(n2529), .config_in(config_chain[7061:7060])); 
mux4 mux_1280 (.in({n2510, n1853, n1830, n592}), .out(n2530), .config_in(config_chain[7063:7062])); 
mux4 mux_1281 (.in({n2551, n1967, n1932, n592}), .out(n2531), .config_in(config_chain[7065:7064])); 
mux4 mux_1282 (.in({n2512, n1855, n1848, n592}), .out(n2532), .config_in(config_chain[7067:7066])); 
mux4 mux_1283 (.in({n2553, n1965, n1934, n592}), .out(n2533), .config_in(config_chain[7069:7068])); 
mux3 mux_1284 (.in({n2514, n1857, n1846}), .out(n2534), .config_in(config_chain[7071:7070])); 
mux3 mux_1285 (.in({n2555, n1963, n1936}), .out(n2535), .config_in(config_chain[7073:7072])); 
mux3 mux_1286 (.in({n2516, n1859, n1844}), .out(n2536), .config_in(config_chain[7075:7074])); 
mux3 mux_1287 (.in({n2557, n1961, n1938}), .out(n2537), .config_in(config_chain[7077:7076])); 
mux3 mux_1288 (.in({n2518, n1861, n1842}), .out(n2538), .config_in(config_chain[7079:7078])); 
mux3 mux_1289 (.in({n2559, n1959, n1940}), .out(n2539), .config_in(config_chain[7081:7080])); 
mux3 mux_1290 (.in({n2520, n1863, n1840}), .out(n2540), .config_in(config_chain[7083:7082])); 
mux3 mux_1291 (.in({n2561, n1957, n1942}), .out(n2541), .config_in(config_chain[7085:7084])); 
mux3 mux_1292 (.in({n2522, n1865, n1838}), .out(n2542), .config_in(config_chain[7087:7086])); 
mux3 mux_1293 (.in({n2563, n1955, n1944}), .out(n2543), .config_in(config_chain[7089:7088])); 
mux3 mux_1294 (.in({n2524, n1867, n1836}), .out(n2544), .config_in(config_chain[7091:7090])); 
mux3 mux_1295 (.in({n2565, n1953, n1946}), .out(n2545), .config_in(config_chain[7093:7092])); 
mux3 mux_1296 (.in({n2526, n1869, n1834}), .out(n2546), .config_in(config_chain[7095:7094])); 
mux3 mux_1297 (.in({n2567, n1951, n1948}), .out(n2547), .config_in(config_chain[7097:7096])); 
mux3 mux_1298 (.in({n2528, n1851, n1832}), .out(n2548), .config_in(config_chain[7099:7098])); 
mux3 mux_1299 (.in({n2569, n1969, n1930}), .out(n2549), .config_in(config_chain[7101:7100])); 
mux4 mux_1300 (.in({n2530, n1953, n1930, n622}), .out(n2550), .config_in(config_chain[7103:7102])); 
mux4 mux_1301 (.in({n2571, n2067, n2032, n622}), .out(n2551), .config_in(config_chain[7105:7104])); 
mux4 mux_1302 (.in({n2532, n1955, n1948, n622}), .out(n2552), .config_in(config_chain[7107:7106])); 
mux4 mux_1303 (.in({n2573, n2065, n2034, n622}), .out(n2553), .config_in(config_chain[7109:7108])); 
mux3 mux_1304 (.in({n2534, n1957, n1946}), .out(n2554), .config_in(config_chain[7111:7110])); 
mux3 mux_1305 (.in({n2575, n2063, n2036}), .out(n2555), .config_in(config_chain[7113:7112])); 
mux3 mux_1306 (.in({n2536, n1959, n1944}), .out(n2556), .config_in(config_chain[7115:7114])); 
mux3 mux_1307 (.in({n2577, n2061, n2038}), .out(n2557), .config_in(config_chain[7117:7116])); 
mux3 mux_1308 (.in({n2538, n1961, n1942}), .out(n2558), .config_in(config_chain[7119:7118])); 
mux3 mux_1309 (.in({n2579, n2059, n2040}), .out(n2559), .config_in(config_chain[7121:7120])); 
mux3 mux_1310 (.in({n2540, n1963, n1940}), .out(n2560), .config_in(config_chain[7123:7122])); 
mux3 mux_1311 (.in({n2581, n2057, n2042}), .out(n2561), .config_in(config_chain[7125:7124])); 
mux3 mux_1312 (.in({n2542, n1965, n1938}), .out(n2562), .config_in(config_chain[7127:7126])); 
mux3 mux_1313 (.in({n2583, n2055, n2044}), .out(n2563), .config_in(config_chain[7129:7128])); 
mux3 mux_1314 (.in({n2544, n1967, n1936}), .out(n2564), .config_in(config_chain[7131:7130])); 
mux3 mux_1315 (.in({n2585, n2053, n2046}), .out(n2565), .config_in(config_chain[7133:7132])); 
mux3 mux_1316 (.in({n2546, n1969, n1934}), .out(n2566), .config_in(config_chain[7135:7134])); 
mux3 mux_1317 (.in({n2587, n2051, n2048}), .out(n2567), .config_in(config_chain[7137:7136])); 
mux3 mux_1318 (.in({n2548, n1951, n1932}), .out(n2568), .config_in(config_chain[7139:7138])); 
mux3 mux_1319 (.in({n2589, n2069, n2030}), .out(n2569), .config_in(config_chain[7141:7140])); 
mux4 mux_1320 (.in({n2550, n2053, n2030, n652}), .out(n2570), .config_in(config_chain[7143:7142])); 
mux4 mux_1321 (.in({n2591, n2167, n2132, n652}), .out(n2571), .config_in(config_chain[7145:7144])); 
mux4 mux_1322 (.in({n2552, n2055, n2048, n652}), .out(n2572), .config_in(config_chain[7147:7146])); 
mux4 mux_1323 (.in({n2593, n2165, n2134, n652}), .out(n2573), .config_in(config_chain[7149:7148])); 
mux3 mux_1324 (.in({n2554, n2057, n2046}), .out(n2574), .config_in(config_chain[7151:7150])); 
mux3 mux_1325 (.in({n2595, n2163, n2136}), .out(n2575), .config_in(config_chain[7153:7152])); 
mux3 mux_1326 (.in({n2556, n2059, n2044}), .out(n2576), .config_in(config_chain[7155:7154])); 
mux3 mux_1327 (.in({n2597, n2161, n2138}), .out(n2577), .config_in(config_chain[7157:7156])); 
mux3 mux_1328 (.in({n2558, n2061, n2042}), .out(n2578), .config_in(config_chain[7159:7158])); 
mux3 mux_1329 (.in({n2599, n2159, n2140}), .out(n2579), .config_in(config_chain[7161:7160])); 
mux3 mux_1330 (.in({n2560, n2063, n2040}), .out(n2580), .config_in(config_chain[7163:7162])); 
mux3 mux_1331 (.in({n2601, n2157, n2142}), .out(n2581), .config_in(config_chain[7165:7164])); 
mux3 mux_1332 (.in({n2562, n2065, n2038}), .out(n2582), .config_in(config_chain[7167:7166])); 
mux3 mux_1333 (.in({n2603, n2155, n2144}), .out(n2583), .config_in(config_chain[7169:7168])); 
mux3 mux_1334 (.in({n2564, n2067, n2036}), .out(n2584), .config_in(config_chain[7171:7170])); 
mux3 mux_1335 (.in({n2605, n2153, n2146}), .out(n2585), .config_in(config_chain[7173:7172])); 
mux3 mux_1336 (.in({n2566, n2069, n2034}), .out(n2586), .config_in(config_chain[7175:7174])); 
mux3 mux_1337 (.in({n2607, n2151, n2148}), .out(n2587), .config_in(config_chain[7177:7176])); 
mux3 mux_1338 (.in({n2568, n2051, n2032}), .out(n2588), .config_in(config_chain[7179:7178])); 
mux3 mux_1339 (.in({n2609, n2169, n2130}), .out(n2589), .config_in(config_chain[7181:7180])); 
mux4 mux_1340 (.in({n2570, n2153, n2130, n682}), .out(n2590), .config_in(config_chain[7183:7182])); 
mux3 mux_1341 (.in({n2251, n2230, n682}), .out(n2591), .config_in(config_chain[7185:7184])); 
mux4 mux_1342 (.in({n2572, n2155, n2148, n682}), .out(n2592), .config_in(config_chain[7187:7186])); 
mux3 mux_1343 (.in({n2259, n2238, n682}), .out(n2593), .config_in(config_chain[7189:7188])); 
mux3 mux_1344 (.in({n2574, n2157, n2146}), .out(n2594), .config_in(config_chain[7191:7190])); 
mux2 mux_1345 (.in({n2261, n2240}), .out(n2595), .config_in(config_chain[7192:7192])); 
mux3 mux_1346 (.in({n2576, n2159, n2144}), .out(n2596), .config_in(config_chain[7194:7193])); 
mux2 mux_1347 (.in({n2253, n2232}), .out(n2597), .config_in(config_chain[7195:7195])); 
mux3 mux_1348 (.in({n2578, n2161, n2142}), .out(n2598), .config_in(config_chain[7197:7196])); 
mux2 mux_1349 (.in({n2263, n2242}), .out(n2599), .config_in(config_chain[7198:7198])); 
mux3 mux_1350 (.in({n2580, n2163, n2140}), .out(n2600), .config_in(config_chain[7200:7199])); 
mux2 mux_1351 (.in({n2265, n2244}), .out(n2601), .config_in(config_chain[7201:7201])); 
mux3 mux_1352 (.in({n2582, n2165, n2138}), .out(n2602), .config_in(config_chain[7203:7202])); 
mux2 mux_1353 (.in({n2255, n2234}), .out(n2603), .config_in(config_chain[7204:7204])); 
mux3 mux_1354 (.in({n2584, n2167, n2136}), .out(n2604), .config_in(config_chain[7206:7205])); 
mux2 mux_1355 (.in({n2267, n2246}), .out(n2605), .config_in(config_chain[7207:7207])); 
mux3 mux_1356 (.in({n2586, n2169, n2134}), .out(n2606), .config_in(config_chain[7209:7208])); 
mux2 mux_1357 (.in({n2269, n2248}), .out(n2607), .config_in(config_chain[7210:7210])); 
mux3 mux_1358 (.in({n2588, n2151, n2132}), .out(n2608), .config_in(config_chain[7212:7211])); 
mux2 mux_1359 (.in({n2257, n2236}), .out(n2609), .config_in(config_chain[7213:7213])); 
mux3 mux_1360 (.in({n1777, n1756, n808}), .out(n2610), .config_in(config_chain[7215:7214])); 
mux4 mux_1361 (.in({n2631, n1887, n1852, n808}), .out(n2611), .config_in(config_chain[7217:7216])); 
mux3 mux_1362 (.in({n1779, n1758, n808}), .out(n2612), .config_in(config_chain[7219:7218])); 
mux4 mux_1363 (.in({n2633, n1885, n1854, n808}), .out(n2613), .config_in(config_chain[7221:7220])); 
mux2 mux_1364 (.in({n1771, n1750}), .out(n2614), .config_in(config_chain[7222:7222])); 
mux3 mux_1365 (.in({n2635, n1883, n1856}), .out(n2615), .config_in(config_chain[7224:7223])); 
mux2 mux_1366 (.in({n1781, n1760}), .out(n2616), .config_in(config_chain[7225:7225])); 
mux3 mux_1367 (.in({n2637, n1881, n1858}), .out(n2617), .config_in(config_chain[7227:7226])); 
mux2 mux_1368 (.in({n1783, n1762}), .out(n2618), .config_in(config_chain[7228:7228])); 
mux3 mux_1369 (.in({n2639, n1879, n1860}), .out(n2619), .config_in(config_chain[7230:7229])); 
mux2 mux_1370 (.in({n1773, n1752}), .out(n2620), .config_in(config_chain[7231:7231])); 
mux3 mux_1371 (.in({n2641, n1877, n1862}), .out(n2621), .config_in(config_chain[7233:7232])); 
mux2 mux_1372 (.in({n1785, n1764}), .out(n2622), .config_in(config_chain[7234:7234])); 
mux3 mux_1373 (.in({n2643, n1875, n1864}), .out(n2623), .config_in(config_chain[7236:7235])); 
mux2 mux_1374 (.in({n1787, n1766}), .out(n2624), .config_in(config_chain[7237:7237])); 
mux3 mux_1375 (.in({n2645, n1873, n1866}), .out(n2625), .config_in(config_chain[7239:7238])); 
mux2 mux_1376 (.in({n1775, n1754}), .out(n2626), .config_in(config_chain[7240:7240])); 
mux3 mux_1377 (.in({n2647, n1871, n1868}), .out(n2627), .config_in(config_chain[7242:7241])); 
mux2 mux_1378 (.in({n1789, n1768}), .out(n2628), .config_in(config_chain[7243:7243])); 
mux3 mux_1379 (.in({n2649, n1889, n1850}), .out(n2629), .config_in(config_chain[7245:7244])); 
mux4 mux_1380 (.in({n2610, n1873, n1850, n838}), .out(n2630), .config_in(config_chain[7247:7246])); 
mux4 mux_1381 (.in({n2651, n1987, n1952, n838}), .out(n2631), .config_in(config_chain[7249:7248])); 
mux4 mux_1382 (.in({n2612, n1875, n1868, n838}), .out(n2632), .config_in(config_chain[7251:7250])); 
mux4 mux_1383 (.in({n2653, n1985, n1954, n838}), .out(n2633), .config_in(config_chain[7253:7252])); 
mux3 mux_1384 (.in({n2614, n1877, n1866}), .out(n2634), .config_in(config_chain[7255:7254])); 
mux3 mux_1385 (.in({n2655, n1983, n1956}), .out(n2635), .config_in(config_chain[7257:7256])); 
mux3 mux_1386 (.in({n2616, n1879, n1864}), .out(n2636), .config_in(config_chain[7259:7258])); 
mux3 mux_1387 (.in({n2657, n1981, n1958}), .out(n2637), .config_in(config_chain[7261:7260])); 
mux3 mux_1388 (.in({n2618, n1881, n1862}), .out(n2638), .config_in(config_chain[7263:7262])); 
mux3 mux_1389 (.in({n2659, n1979, n1960}), .out(n2639), .config_in(config_chain[7265:7264])); 
mux3 mux_1390 (.in({n2620, n1883, n1860}), .out(n2640), .config_in(config_chain[7267:7266])); 
mux3 mux_1391 (.in({n2661, n1977, n1962}), .out(n2641), .config_in(config_chain[7269:7268])); 
mux3 mux_1392 (.in({n2622, n1885, n1858}), .out(n2642), .config_in(config_chain[7271:7270])); 
mux3 mux_1393 (.in({n2663, n1975, n1964}), .out(n2643), .config_in(config_chain[7273:7272])); 
mux3 mux_1394 (.in({n2624, n1887, n1856}), .out(n2644), .config_in(config_chain[7275:7274])); 
mux3 mux_1395 (.in({n2665, n1973, n1966}), .out(n2645), .config_in(config_chain[7277:7276])); 
mux3 mux_1396 (.in({n2626, n1889, n1854}), .out(n2646), .config_in(config_chain[7279:7278])); 
mux3 mux_1397 (.in({n2667, n1971, n1968}), .out(n2647), .config_in(config_chain[7281:7280])); 
mux3 mux_1398 (.in({n2628, n1871, n1852}), .out(n2648), .config_in(config_chain[7283:7282])); 
mux3 mux_1399 (.in({n2669, n1989, n1950}), .out(n2649), .config_in(config_chain[7285:7284])); 
mux4 mux_1400 (.in({n2630, n1973, n1950, n868}), .out(n2650), .config_in(config_chain[7287:7286])); 
mux4 mux_1401 (.in({n2671, n2087, n2052, n868}), .out(n2651), .config_in(config_chain[7289:7288])); 
mux4 mux_1402 (.in({n2632, n1975, n1968, n868}), .out(n2652), .config_in(config_chain[7291:7290])); 
mux4 mux_1403 (.in({n2673, n2085, n2054, n868}), .out(n2653), .config_in(config_chain[7293:7292])); 
mux3 mux_1404 (.in({n2634, n1977, n1966}), .out(n2654), .config_in(config_chain[7295:7294])); 
mux3 mux_1405 (.in({n2675, n2083, n2056}), .out(n2655), .config_in(config_chain[7297:7296])); 
mux3 mux_1406 (.in({n2636, n1979, n1964}), .out(n2656), .config_in(config_chain[7299:7298])); 
mux3 mux_1407 (.in({n2677, n2081, n2058}), .out(n2657), .config_in(config_chain[7301:7300])); 
mux3 mux_1408 (.in({n2638, n1981, n1962}), .out(n2658), .config_in(config_chain[7303:7302])); 
mux3 mux_1409 (.in({n2679, n2079, n2060}), .out(n2659), .config_in(config_chain[7305:7304])); 
mux3 mux_1410 (.in({n2640, n1983, n1960}), .out(n2660), .config_in(config_chain[7307:7306])); 
mux3 mux_1411 (.in({n2681, n2077, n2062}), .out(n2661), .config_in(config_chain[7309:7308])); 
mux3 mux_1412 (.in({n2642, n1985, n1958}), .out(n2662), .config_in(config_chain[7311:7310])); 
mux3 mux_1413 (.in({n2683, n2075, n2064}), .out(n2663), .config_in(config_chain[7313:7312])); 
mux3 mux_1414 (.in({n2644, n1987, n1956}), .out(n2664), .config_in(config_chain[7315:7314])); 
mux3 mux_1415 (.in({n2685, n2073, n2066}), .out(n2665), .config_in(config_chain[7317:7316])); 
mux3 mux_1416 (.in({n2646, n1989, n1954}), .out(n2666), .config_in(config_chain[7319:7318])); 
mux3 mux_1417 (.in({n2687, n2071, n2068}), .out(n2667), .config_in(config_chain[7321:7320])); 
mux3 mux_1418 (.in({n2648, n1971, n1952}), .out(n2668), .config_in(config_chain[7323:7322])); 
mux3 mux_1419 (.in({n2689, n2089, n2050}), .out(n2669), .config_in(config_chain[7325:7324])); 
mux4 mux_1420 (.in({n2650, n2073, n2050, n898}), .out(n2670), .config_in(config_chain[7327:7326])); 
mux4 mux_1421 (.in({n2691, n2187, n2152, n898}), .out(n2671), .config_in(config_chain[7329:7328])); 
mux4 mux_1422 (.in({n2652, n2075, n2068, n898}), .out(n2672), .config_in(config_chain[7331:7330])); 
mux4 mux_1423 (.in({n2693, n2185, n2154, n898}), .out(n2673), .config_in(config_chain[7333:7332])); 
mux3 mux_1424 (.in({n2654, n2077, n2066}), .out(n2674), .config_in(config_chain[7335:7334])); 
mux3 mux_1425 (.in({n2695, n2183, n2156}), .out(n2675), .config_in(config_chain[7337:7336])); 
mux3 mux_1426 (.in({n2656, n2079, n2064}), .out(n2676), .config_in(config_chain[7339:7338])); 
mux3 mux_1427 (.in({n2697, n2181, n2158}), .out(n2677), .config_in(config_chain[7341:7340])); 
mux3 mux_1428 (.in({n2658, n2081, n2062}), .out(n2678), .config_in(config_chain[7343:7342])); 
mux3 mux_1429 (.in({n2699, n2179, n2160}), .out(n2679), .config_in(config_chain[7345:7344])); 
mux3 mux_1430 (.in({n2660, n2083, n2060}), .out(n2680), .config_in(config_chain[7347:7346])); 
mux3 mux_1431 (.in({n2701, n2177, n2162}), .out(n2681), .config_in(config_chain[7349:7348])); 
mux3 mux_1432 (.in({n2662, n2085, n2058}), .out(n2682), .config_in(config_chain[7351:7350])); 
mux3 mux_1433 (.in({n2703, n2175, n2164}), .out(n2683), .config_in(config_chain[7353:7352])); 
mux3 mux_1434 (.in({n2664, n2087, n2056}), .out(n2684), .config_in(config_chain[7355:7354])); 
mux3 mux_1435 (.in({n2705, n2173, n2166}), .out(n2685), .config_in(config_chain[7357:7356])); 
mux3 mux_1436 (.in({n2666, n2089, n2054}), .out(n2686), .config_in(config_chain[7359:7358])); 
mux3 mux_1437 (.in({n2707, n2171, n2168}), .out(n2687), .config_in(config_chain[7361:7360])); 
mux3 mux_1438 (.in({n2668, n2071, n2052}), .out(n2688), .config_in(config_chain[7363:7362])); 
mux3 mux_1439 (.in({n2709, n2189, n2150}), .out(n2689), .config_in(config_chain[7365:7364])); 
mux4 mux_1440 (.in({n2670, n2173, n2150, n928}), .out(n2690), .config_in(config_chain[7367:7366])); 
mux3 mux_1441 (.in({n2271, n2250, n928}), .out(n2691), .config_in(config_chain[7369:7368])); 
mux4 mux_1442 (.in({n2672, n2175, n2168, n928}), .out(n2692), .config_in(config_chain[7371:7370])); 
mux3 mux_1443 (.in({n2279, n2258, n928}), .out(n2693), .config_in(config_chain[7373:7372])); 
mux3 mux_1444 (.in({n2674, n2177, n2166}), .out(n2694), .config_in(config_chain[7375:7374])); 
mux2 mux_1445 (.in({n2281, n2260}), .out(n2695), .config_in(config_chain[7376:7376])); 
mux3 mux_1446 (.in({n2676, n2179, n2164}), .out(n2696), .config_in(config_chain[7378:7377])); 
mux2 mux_1447 (.in({n2273, n2252}), .out(n2697), .config_in(config_chain[7379:7379])); 
mux3 mux_1448 (.in({n2678, n2181, n2162}), .out(n2698), .config_in(config_chain[7381:7380])); 
mux2 mux_1449 (.in({n2283, n2262}), .out(n2699), .config_in(config_chain[7382:7382])); 
mux3 mux_1450 (.in({n2680, n2183, n2160}), .out(n2700), .config_in(config_chain[7384:7383])); 
mux2 mux_1451 (.in({n2285, n2264}), .out(n2701), .config_in(config_chain[7385:7385])); 
mux3 mux_1452 (.in({n2682, n2185, n2158}), .out(n2702), .config_in(config_chain[7387:7386])); 
mux2 mux_1453 (.in({n2275, n2254}), .out(n2703), .config_in(config_chain[7388:7388])); 
mux3 mux_1454 (.in({n2684, n2187, n2156}), .out(n2704), .config_in(config_chain[7390:7389])); 
mux2 mux_1455 (.in({n2287, n2266}), .out(n2705), .config_in(config_chain[7391:7391])); 
mux3 mux_1456 (.in({n2686, n2189, n2154}), .out(n2706), .config_in(config_chain[7393:7392])); 
mux2 mux_1457 (.in({n2289, n2268}), .out(n2707), .config_in(config_chain[7394:7394])); 
mux3 mux_1458 (.in({n2688, n2171, n2152}), .out(n2708), .config_in(config_chain[7396:7395])); 
mux2 mux_1459 (.in({n2277, n2256}), .out(n2709), .config_in(config_chain[7397:7397])); 
mux3 mux_1460 (.in({n1797, n1776, n1054}), .out(n2710), .config_in(config_chain[7399:7398])); 
mux4 mux_1461 (.in({n2731, n1907, n1872, n1054}), .out(n2711), .config_in(config_chain[7401:7400])); 
mux3 mux_1462 (.in({n1799, n1778, n1054}), .out(n2712), .config_in(config_chain[7403:7402])); 
mux4 mux_1463 (.in({n2733, n1905, n1874, n1054}), .out(n2713), .config_in(config_chain[7405:7404])); 
mux2 mux_1464 (.in({n1791, n1770}), .out(n2714), .config_in(config_chain[7406:7406])); 
mux3 mux_1465 (.in({n2735, n1903, n1876}), .out(n2715), .config_in(config_chain[7408:7407])); 
mux2 mux_1466 (.in({n1801, n1780}), .out(n2716), .config_in(config_chain[7409:7409])); 
mux3 mux_1467 (.in({n2737, n1901, n1878}), .out(n2717), .config_in(config_chain[7411:7410])); 
mux2 mux_1468 (.in({n1803, n1782}), .out(n2718), .config_in(config_chain[7412:7412])); 
mux3 mux_1469 (.in({n2739, n1899, n1880}), .out(n2719), .config_in(config_chain[7414:7413])); 
mux2 mux_1470 (.in({n1793, n1772}), .out(n2720), .config_in(config_chain[7415:7415])); 
mux3 mux_1471 (.in({n2741, n1897, n1882}), .out(n2721), .config_in(config_chain[7417:7416])); 
mux2 mux_1472 (.in({n1805, n1784}), .out(n2722), .config_in(config_chain[7418:7418])); 
mux3 mux_1473 (.in({n2743, n1895, n1884}), .out(n2723), .config_in(config_chain[7420:7419])); 
mux2 mux_1474 (.in({n1807, n1786}), .out(n2724), .config_in(config_chain[7421:7421])); 
mux3 mux_1475 (.in({n2745, n1893, n1886}), .out(n2725), .config_in(config_chain[7423:7422])); 
mux2 mux_1476 (.in({n1795, n1774}), .out(n2726), .config_in(config_chain[7424:7424])); 
mux3 mux_1477 (.in({n2747, n1891, n1888}), .out(n2727), .config_in(config_chain[7426:7425])); 
mux2 mux_1478 (.in({n1809, n1788}), .out(n2728), .config_in(config_chain[7427:7427])); 
mux3 mux_1479 (.in({n2749, n1909, n1870}), .out(n2729), .config_in(config_chain[7429:7428])); 
mux4 mux_1480 (.in({n2710, n1893, n1870, n1084}), .out(n2730), .config_in(config_chain[7431:7430])); 
mux4 mux_1481 (.in({n2751, n2007, n1972, n1084}), .out(n2731), .config_in(config_chain[7433:7432])); 
mux4 mux_1482 (.in({n2712, n1895, n1888, n1084}), .out(n2732), .config_in(config_chain[7435:7434])); 
mux4 mux_1483 (.in({n2753, n2005, n1974, n1084}), .out(n2733), .config_in(config_chain[7437:7436])); 
mux3 mux_1484 (.in({n2714, n1897, n1886}), .out(n2734), .config_in(config_chain[7439:7438])); 
mux3 mux_1485 (.in({n2755, n2003, n1976}), .out(n2735), .config_in(config_chain[7441:7440])); 
mux3 mux_1486 (.in({n2716, n1899, n1884}), .out(n2736), .config_in(config_chain[7443:7442])); 
mux3 mux_1487 (.in({n2757, n2001, n1978}), .out(n2737), .config_in(config_chain[7445:7444])); 
mux3 mux_1488 (.in({n2718, n1901, n1882}), .out(n2738), .config_in(config_chain[7447:7446])); 
mux3 mux_1489 (.in({n2759, n1999, n1980}), .out(n2739), .config_in(config_chain[7449:7448])); 
mux3 mux_1490 (.in({n2720, n1903, n1880}), .out(n2740), .config_in(config_chain[7451:7450])); 
mux3 mux_1491 (.in({n2761, n1997, n1982}), .out(n2741), .config_in(config_chain[7453:7452])); 
mux3 mux_1492 (.in({n2722, n1905, n1878}), .out(n2742), .config_in(config_chain[7455:7454])); 
mux3 mux_1493 (.in({n2763, n1995, n1984}), .out(n2743), .config_in(config_chain[7457:7456])); 
mux3 mux_1494 (.in({n2724, n1907, n1876}), .out(n2744), .config_in(config_chain[7459:7458])); 
mux3 mux_1495 (.in({n2765, n1993, n1986}), .out(n2745), .config_in(config_chain[7461:7460])); 
mux3 mux_1496 (.in({n2726, n1909, n1874}), .out(n2746), .config_in(config_chain[7463:7462])); 
mux3 mux_1497 (.in({n2767, n1991, n1988}), .out(n2747), .config_in(config_chain[7465:7464])); 
mux3 mux_1498 (.in({n2728, n1891, n1872}), .out(n2748), .config_in(config_chain[7467:7466])); 
mux3 mux_1499 (.in({n2769, n2009, n1970}), .out(n2749), .config_in(config_chain[7469:7468])); 
mux4 mux_1500 (.in({n2730, n1993, n1970, n1114}), .out(n2750), .config_in(config_chain[7471:7470])); 
mux4 mux_1501 (.in({n2771, n2107, n2072, n1114}), .out(n2751), .config_in(config_chain[7473:7472])); 
mux4 mux_1502 (.in({n2732, n1995, n1988, n1114}), .out(n2752), .config_in(config_chain[7475:7474])); 
mux4 mux_1503 (.in({n2773, n2105, n2074, n1114}), .out(n2753), .config_in(config_chain[7477:7476])); 
mux3 mux_1504 (.in({n2734, n1997, n1986}), .out(n2754), .config_in(config_chain[7479:7478])); 
mux3 mux_1505 (.in({n2775, n2103, n2076}), .out(n2755), .config_in(config_chain[7481:7480])); 
mux3 mux_1506 (.in({n2736, n1999, n1984}), .out(n2756), .config_in(config_chain[7483:7482])); 
mux3 mux_1507 (.in({n2777, n2101, n2078}), .out(n2757), .config_in(config_chain[7485:7484])); 
mux3 mux_1508 (.in({n2738, n2001, n1982}), .out(n2758), .config_in(config_chain[7487:7486])); 
mux3 mux_1509 (.in({n2779, n2099, n2080}), .out(n2759), .config_in(config_chain[7489:7488])); 
mux3 mux_1510 (.in({n2740, n2003, n1980}), .out(n2760), .config_in(config_chain[7491:7490])); 
mux3 mux_1511 (.in({n2781, n2097, n2082}), .out(n2761), .config_in(config_chain[7493:7492])); 
mux3 mux_1512 (.in({n2742, n2005, n1978}), .out(n2762), .config_in(config_chain[7495:7494])); 
mux3 mux_1513 (.in({n2783, n2095, n2084}), .out(n2763), .config_in(config_chain[7497:7496])); 
mux3 mux_1514 (.in({n2744, n2007, n1976}), .out(n2764), .config_in(config_chain[7499:7498])); 
mux3 mux_1515 (.in({n2785, n2093, n2086}), .out(n2765), .config_in(config_chain[7501:7500])); 
mux3 mux_1516 (.in({n2746, n2009, n1974}), .out(n2766), .config_in(config_chain[7503:7502])); 
mux3 mux_1517 (.in({n2787, n2091, n2088}), .out(n2767), .config_in(config_chain[7505:7504])); 
mux3 mux_1518 (.in({n2748, n1991, n1972}), .out(n2768), .config_in(config_chain[7507:7506])); 
mux3 mux_1519 (.in({n2789, n2109, n2070}), .out(n2769), .config_in(config_chain[7509:7508])); 
mux4 mux_1520 (.in({n2750, n2093, n2070, n1144}), .out(n2770), .config_in(config_chain[7511:7510])); 
mux4 mux_1521 (.in({n2791, n2207, n2172, n1144}), .out(n2771), .config_in(config_chain[7513:7512])); 
mux4 mux_1522 (.in({n2752, n2095, n2088, n1144}), .out(n2772), .config_in(config_chain[7515:7514])); 
mux4 mux_1523 (.in({n2793, n2205, n2174, n1144}), .out(n2773), .config_in(config_chain[7517:7516])); 
mux3 mux_1524 (.in({n2754, n2097, n2086}), .out(n2774), .config_in(config_chain[7519:7518])); 
mux3 mux_1525 (.in({n2795, n2203, n2176}), .out(n2775), .config_in(config_chain[7521:7520])); 
mux3 mux_1526 (.in({n2756, n2099, n2084}), .out(n2776), .config_in(config_chain[7523:7522])); 
mux3 mux_1527 (.in({n2797, n2201, n2178}), .out(n2777), .config_in(config_chain[7525:7524])); 
mux3 mux_1528 (.in({n2758, n2101, n2082}), .out(n2778), .config_in(config_chain[7527:7526])); 
mux3 mux_1529 (.in({n2799, n2199, n2180}), .out(n2779), .config_in(config_chain[7529:7528])); 
mux3 mux_1530 (.in({n2760, n2103, n2080}), .out(n2780), .config_in(config_chain[7531:7530])); 
mux3 mux_1531 (.in({n2801, n2197, n2182}), .out(n2781), .config_in(config_chain[7533:7532])); 
mux3 mux_1532 (.in({n2762, n2105, n2078}), .out(n2782), .config_in(config_chain[7535:7534])); 
mux3 mux_1533 (.in({n2803, n2195, n2184}), .out(n2783), .config_in(config_chain[7537:7536])); 
mux3 mux_1534 (.in({n2764, n2107, n2076}), .out(n2784), .config_in(config_chain[7539:7538])); 
mux3 mux_1535 (.in({n2805, n2193, n2186}), .out(n2785), .config_in(config_chain[7541:7540])); 
mux3 mux_1536 (.in({n2766, n2109, n2074}), .out(n2786), .config_in(config_chain[7543:7542])); 
mux3 mux_1537 (.in({n2807, n2191, n2188}), .out(n2787), .config_in(config_chain[7545:7544])); 
mux3 mux_1538 (.in({n2768, n2091, n2072}), .out(n2788), .config_in(config_chain[7547:7546])); 
mux3 mux_1539 (.in({n2809, n2209, n2170}), .out(n2789), .config_in(config_chain[7549:7548])); 
mux4 mux_1540 (.in({n2770, n2193, n2170, n1174}), .out(n2790), .config_in(config_chain[7551:7550])); 
mux3 mux_1541 (.in({n2291, n2270, n1174}), .out(n2791), .config_in(config_chain[7553:7552])); 
mux4 mux_1542 (.in({n2772, n2195, n2188, n1174}), .out(n2792), .config_in(config_chain[7555:7554])); 
mux3 mux_1543 (.in({n2299, n2278, n1174}), .out(n2793), .config_in(config_chain[7557:7556])); 
mux3 mux_1544 (.in({n2774, n2197, n2186}), .out(n2794), .config_in(config_chain[7559:7558])); 
mux2 mux_1545 (.in({n2301, n2280}), .out(n2795), .config_in(config_chain[7560:7560])); 
mux3 mux_1546 (.in({n2776, n2199, n2184}), .out(n2796), .config_in(config_chain[7562:7561])); 
mux2 mux_1547 (.in({n2293, n2272}), .out(n2797), .config_in(config_chain[7563:7563])); 
mux3 mux_1548 (.in({n2778, n2201, n2182}), .out(n2798), .config_in(config_chain[7565:7564])); 
mux2 mux_1549 (.in({n2303, n2282}), .out(n2799), .config_in(config_chain[7566:7566])); 
mux3 mux_1550 (.in({n2780, n2203, n2180}), .out(n2800), .config_in(config_chain[7568:7567])); 
mux2 mux_1551 (.in({n2305, n2284}), .out(n2801), .config_in(config_chain[7569:7569])); 
mux3 mux_1552 (.in({n2782, n2205, n2178}), .out(n2802), .config_in(config_chain[7571:7570])); 
mux2 mux_1553 (.in({n2295, n2274}), .out(n2803), .config_in(config_chain[7572:7572])); 
mux3 mux_1554 (.in({n2784, n2207, n2176}), .out(n2804), .config_in(config_chain[7574:7573])); 
mux2 mux_1555 (.in({n2307, n2286}), .out(n2805), .config_in(config_chain[7575:7575])); 
mux3 mux_1556 (.in({n2786, n2209, n2174}), .out(n2806), .config_in(config_chain[7577:7576])); 
mux2 mux_1557 (.in({n2309, n2288}), .out(n2807), .config_in(config_chain[7578:7578])); 
mux3 mux_1558 (.in({n2788, n2191, n2172}), .out(n2808), .config_in(config_chain[7580:7579])); 
mux2 mux_1559 (.in({n2297, n2276}), .out(n2809), .config_in(config_chain[7581:7581])); 
mux3 mux_1560 (.in({n1790, n1507, n1300}), .out(n2810), .config_in(config_chain[7583:7582])); 
mux4 mux_1561 (.in({n2831, n1890, n1507, n1300}), .out(n2811), .config_in(config_chain[7585:7584])); 
mux3 mux_1562 (.in({n1808, n1507, n1300}), .out(n2812), .config_in(config_chain[7587:7586])); 
mux4 mux_1563 (.in({n2833, n1892, n1507, n1300}), .out(n2813), .config_in(config_chain[7589:7588])); 
mux3 mux_1564 (.in({n1806, n1510, n1495}), .out(n2814), .config_in(config_chain[7591:7590])); 
mux4 mux_1565 (.in({n2835, n1894, n1510, n1495}), .out(n2815), .config_in(config_chain[7593:7592])); 
mux3 mux_1566 (.in({n1804, n1510, n1495}), .out(n2816), .config_in(config_chain[7595:7594])); 
mux4 mux_1567 (.in({n2837, n1896, n1510, n1495}), .out(n2817), .config_in(config_chain[7597:7596])); 
mux3 mux_1568 (.in({n1802, n1513, n1498}), .out(n2818), .config_in(config_chain[7599:7598])); 
mux4 mux_1569 (.in({n2839, n1898, n1513, n1498}), .out(n2819), .config_in(config_chain[7601:7600])); 
mux3 mux_1570 (.in({n1800, n1513, n1498}), .out(n2820), .config_in(config_chain[7603:7602])); 
mux4 mux_1571 (.in({n2841, n1900, n1513, n1498}), .out(n2821), .config_in(config_chain[7605:7604])); 
mux3 mux_1572 (.in({n1798, n1516, n1501}), .out(n2822), .config_in(config_chain[7607:7606])); 
mux4 mux_1573 (.in({n2843, n1902, n1516, n1501}), .out(n2823), .config_in(config_chain[7609:7608])); 
mux3 mux_1574 (.in({n1796, n1516, n1501}), .out(n2824), .config_in(config_chain[7611:7610])); 
mux4 mux_1575 (.in({n2845, n1904, n1516, n1501}), .out(n2825), .config_in(config_chain[7613:7612])); 
mux2 mux_1576 (.in({n1794, n1504}), .out(n2826), .config_in(config_chain[7614:7614])); 
mux3 mux_1577 (.in({n2847, n1906, n1504}), .out(n2827), .config_in(config_chain[7616:7615])); 
mux2 mux_1578 (.in({n1792, n1504}), .out(n2828), .config_in(config_chain[7617:7617])); 
mux3 mux_1579 (.in({n2849, n1908, n1504}), .out(n2829), .config_in(config_chain[7619:7618])); 
mux4 mux_1580 (.in({n2810, n1890, n1555, n1330}), .out(n2830), .config_in(config_chain[7621:7620])); 
mux4 mux_1581 (.in({n2851, n1990, n1555, n1330}), .out(n2831), .config_in(config_chain[7623:7622])); 
mux4 mux_1582 (.in({n2812, n1892, n1555, n1330}), .out(n2832), .config_in(config_chain[7625:7624])); 
mux4 mux_1583 (.in({n2853, n1992, n1555, n1330}), .out(n2833), .config_in(config_chain[7627:7626])); 
mux4 mux_1584 (.in({n2814, n1894, n1558, n1543}), .out(n2834), .config_in(config_chain[7629:7628])); 
mux4 mux_1585 (.in({n2855, n1994, n1558, n1543}), .out(n2835), .config_in(config_chain[7631:7630])); 
mux4 mux_1586 (.in({n2816, n1896, n1558, n1543}), .out(n2836), .config_in(config_chain[7633:7632])); 
mux4 mux_1587 (.in({n2857, n1996, n1558, n1543}), .out(n2837), .config_in(config_chain[7635:7634])); 
mux4 mux_1588 (.in({n2818, n1898, n1561, n1546}), .out(n2838), .config_in(config_chain[7637:7636])); 
mux4 mux_1589 (.in({n2859, n1998, n1561, n1546}), .out(n2839), .config_in(config_chain[7639:7638])); 
mux4 mux_1590 (.in({n2820, n1900, n1561, n1546}), .out(n2840), .config_in(config_chain[7641:7640])); 
mux4 mux_1591 (.in({n2861, n2000, n1561, n1546}), .out(n2841), .config_in(config_chain[7643:7642])); 
mux4 mux_1592 (.in({n2822, n1902, n1564, n1549}), .out(n2842), .config_in(config_chain[7645:7644])); 
mux4 mux_1593 (.in({n2863, n2002, n1564, n1549}), .out(n2843), .config_in(config_chain[7647:7646])); 
mux4 mux_1594 (.in({n2824, n1904, n1564, n1549}), .out(n2844), .config_in(config_chain[7649:7648])); 
mux4 mux_1595 (.in({n2865, n2004, n1564, n1549}), .out(n2845), .config_in(config_chain[7651:7650])); 
mux3 mux_1596 (.in({n2826, n1906, n1552}), .out(n2846), .config_in(config_chain[7653:7652])); 
mux3 mux_1597 (.in({n2867, n2006, n1552}), .out(n2847), .config_in(config_chain[7655:7654])); 
mux3 mux_1598 (.in({n2828, n1908, n1552}), .out(n2848), .config_in(config_chain[7657:7656])); 
mux3 mux_1599 (.in({n2869, n2008, n1552}), .out(n2849), .config_in(config_chain[7659:7658])); 
mux4 mux_1600 (.in({n2830, n1990, n1603, n1360}), .out(n2850), .config_in(config_chain[7661:7660])); 
mux4 mux_1601 (.in({n2871, n2090, n1603, n1360}), .out(n2851), .config_in(config_chain[7663:7662])); 
mux4 mux_1602 (.in({n2832, n1992, n1603, n1360}), .out(n2852), .config_in(config_chain[7665:7664])); 
mux4 mux_1603 (.in({n2873, n2092, n1603, n1360}), .out(n2853), .config_in(config_chain[7667:7666])); 
mux4 mux_1604 (.in({n2834, n1994, n1606, n1591}), .out(n2854), .config_in(config_chain[7669:7668])); 
mux4 mux_1605 (.in({n2875, n2094, n1606, n1591}), .out(n2855), .config_in(config_chain[7671:7670])); 
mux4 mux_1606 (.in({n2836, n1996, n1606, n1591}), .out(n2856), .config_in(config_chain[7673:7672])); 
mux4 mux_1607 (.in({n2877, n2096, n1606, n1591}), .out(n2857), .config_in(config_chain[7675:7674])); 
mux4 mux_1608 (.in({n2838, n1998, n1609, n1594}), .out(n2858), .config_in(config_chain[7677:7676])); 
mux4 mux_1609 (.in({n2879, n2098, n1609, n1594}), .out(n2859), .config_in(config_chain[7679:7678])); 
mux4 mux_1610 (.in({n2840, n2000, n1609, n1594}), .out(n2860), .config_in(config_chain[7681:7680])); 
mux4 mux_1611 (.in({n2881, n2100, n1609, n1594}), .out(n2861), .config_in(config_chain[7683:7682])); 
mux4 mux_1612 (.in({n2842, n2002, n1612, n1597}), .out(n2862), .config_in(config_chain[7685:7684])); 
mux4 mux_1613 (.in({n2883, n2102, n1612, n1597}), .out(n2863), .config_in(config_chain[7687:7686])); 
mux4 mux_1614 (.in({n2844, n2004, n1612, n1597}), .out(n2864), .config_in(config_chain[7689:7688])); 
mux4 mux_1615 (.in({n2885, n2104, n1612, n1597}), .out(n2865), .config_in(config_chain[7691:7690])); 
mux3 mux_1616 (.in({n2846, n2006, n1600}), .out(n2866), .config_in(config_chain[7693:7692])); 
mux3 mux_1617 (.in({n2887, n2106, n1600}), .out(n2867), .config_in(config_chain[7695:7694])); 
mux3 mux_1618 (.in({n2848, n2008, n1600}), .out(n2868), .config_in(config_chain[7697:7696])); 
mux3 mux_1619 (.in({n2889, n2108, n1600}), .out(n2869), .config_in(config_chain[7699:7698])); 
mux4 mux_1620 (.in({n2850, n2090, n1651, n1390}), .out(n2870), .config_in(config_chain[7701:7700])); 
mux4 mux_1621 (.in({n2891, n2190, n1651, n1390}), .out(n2871), .config_in(config_chain[7703:7702])); 
mux4 mux_1622 (.in({n2852, n2092, n1651, n1390}), .out(n2872), .config_in(config_chain[7705:7704])); 
mux4 mux_1623 (.in({n2893, n2192, n1651, n1390}), .out(n2873), .config_in(config_chain[7707:7706])); 
mux4 mux_1624 (.in({n2854, n2094, n1654, n1639}), .out(n2874), .config_in(config_chain[7709:7708])); 
mux4 mux_1625 (.in({n2895, n2194, n1654, n1639}), .out(n2875), .config_in(config_chain[7711:7710])); 
mux4 mux_1626 (.in({n2856, n2096, n1654, n1639}), .out(n2876), .config_in(config_chain[7713:7712])); 
mux4 mux_1627 (.in({n2897, n2196, n1654, n1639}), .out(n2877), .config_in(config_chain[7715:7714])); 
mux4 mux_1628 (.in({n2858, n2098, n1657, n1642}), .out(n2878), .config_in(config_chain[7717:7716])); 
mux4 mux_1629 (.in({n2899, n2198, n1657, n1642}), .out(n2879), .config_in(config_chain[7719:7718])); 
mux4 mux_1630 (.in({n2860, n2100, n1657, n1642}), .out(n2880), .config_in(config_chain[7721:7720])); 
mux4 mux_1631 (.in({n2901, n2200, n1657, n1642}), .out(n2881), .config_in(config_chain[7723:7722])); 
mux4 mux_1632 (.in({n2862, n2102, n1660, n1645}), .out(n2882), .config_in(config_chain[7725:7724])); 
mux4 mux_1633 (.in({n2903, n2202, n1660, n1645}), .out(n2883), .config_in(config_chain[7727:7726])); 
mux4 mux_1634 (.in({n2864, n2104, n1660, n1645}), .out(n2884), .config_in(config_chain[7729:7728])); 
mux4 mux_1635 (.in({n2905, n2204, n1660, n1645}), .out(n2885), .config_in(config_chain[7731:7730])); 
mux3 mux_1636 (.in({n2866, n2106, n1648}), .out(n2886), .config_in(config_chain[7733:7732])); 
mux3 mux_1637 (.in({n2907, n2206, n1648}), .out(n2887), .config_in(config_chain[7735:7734])); 
mux3 mux_1638 (.in({n2868, n2108, n1648}), .out(n2888), .config_in(config_chain[7737:7736])); 
mux3 mux_1639 (.in({n2909, n2208, n1648}), .out(n2889), .config_in(config_chain[7739:7738])); 
mux4 mux_1640 (.in({n2870, n2190, n1699, n1420}), .out(n2890), .config_in(config_chain[7741:7740])); 
mux3 mux_1641 (.in({n2292, n1699, n1420}), .out(n2891), .config_in(config_chain[7743:7742])); 
mux4 mux_1642 (.in({n2872, n2192, n1699, n1420}), .out(n2892), .config_in(config_chain[7745:7744])); 
mux3 mux_1643 (.in({n2294, n1699, n1420}), .out(n2893), .config_in(config_chain[7747:7746])); 
mux4 mux_1644 (.in({n2874, n2194, n1702, n1687}), .out(n2894), .config_in(config_chain[7749:7748])); 
mux3 mux_1645 (.in({n2296, n1702, n1687}), .out(n2895), .config_in(config_chain[7751:7750])); 
mux4 mux_1646 (.in({n2876, n2196, n1702, n1687}), .out(n2896), .config_in(config_chain[7753:7752])); 
mux3 mux_1647 (.in({n2298, n1702, n1687}), .out(n2897), .config_in(config_chain[7755:7754])); 
mux4 mux_1648 (.in({n2878, n2198, n1705, n1690}), .out(n2898), .config_in(config_chain[7757:7756])); 
mux3 mux_1649 (.in({n2300, n1705, n1690}), .out(n2899), .config_in(config_chain[7759:7758])); 
mux4 mux_1650 (.in({n2880, n2200, n1705, n1690}), .out(n2900), .config_in(config_chain[7761:7760])); 
mux3 mux_1651 (.in({n2302, n1705, n1690}), .out(n2901), .config_in(config_chain[7763:7762])); 
mux4 mux_1652 (.in({n2882, n2202, n1708, n1693}), .out(n2902), .config_in(config_chain[7765:7764])); 
mux3 mux_1653 (.in({n2304, n1708, n1693}), .out(n2903), .config_in(config_chain[7767:7766])); 
mux4 mux_1654 (.in({n2884, n2204, n1708, n1693}), .out(n2904), .config_in(config_chain[7769:7768])); 
mux3 mux_1655 (.in({n2306, n1708, n1693}), .out(n2905), .config_in(config_chain[7771:7770])); 
mux3 mux_1656 (.in({n2886, n2206, n1696}), .out(n2906), .config_in(config_chain[7773:7772])); 
mux2 mux_1657 (.in({n2308, n1696}), .out(n2907), .config_in(config_chain[7774:7774])); 
mux3 mux_1658 (.in({n2888, n2208, n1696}), .out(n2908), .config_in(config_chain[7776:7775])); 
mux2 mux_1659 (.in({n2290, n1696}), .out(n2909), .config_in(config_chain[7777:7777])); 

wire [7777:0]config_chain_shift;
assign config_chain = config_en?0:config_chain_shift;
config_helper config_helper_0 ( .config_in(config_in), .config_out(config_chain_shift[7777:0]), .config_en(config_en), .reset(reset), .clk(config_clk) );

endmodule

module config_helper (
	input clk,
	input reset,
	input config_in,
	input config_en,
	output [7777:0]config_out
);

latch config_latch_start ( .clk(clk), .reset(reset), .en(config_en), .in(config_in), .out(config_out[0]) );
generate
genvar i;
for(i=0; i<7778; i=i+2)
begin: shifter1
latch config_latch ( .clk(clk), .reset(reset), .en(config_en), .in(config_out[i]), .out(config_out[i+1]) );
end
endgenerate

generate
for(i=1; i<7777; i=i+2)
begin: shifter2
latch config_latch ( .clk(clk), .reset(reset), .en(config_en), .in(config_out[i]), .out(config_out[i+1]) );
end
endgenerate

endmodule
